module forward_jump(
	
);
//input output
	input EXMEM_RegWrite;
	input EXMEM_Reg
//reg & wire
//combinatinal
//no sequentioal
endmodule
