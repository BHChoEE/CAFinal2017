module Control();
end module
