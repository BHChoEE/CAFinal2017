
module Control ( inst, funct, eq, PCSrc, IF_Flush, RegWrite, ALURsc, ALUOp, 
        RegDst, MemWrite, MemRead, MemtoReg, Jump, JumpR, raWrite, Branch, 
        Shift, Mul, Div, HI, LO );
  input [5:0] inst;
  input [5:0] funct;
  output [1:0] ALUOp;
  input eq;
  output PCSrc, IF_Flush, RegWrite, ALURsc, RegDst, MemWrite, MemRead,
         MemtoReg, Jump, JumpR, raWrite, Branch, Shift, Mul, Div, HI, LO;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n5, n6, n7, n8, n9, n32, n33,
         n34, n35;

  CLKINVX1 U3 ( .A(inst[2]), .Y(n32) );
  NAND4X1 U4 ( .A(funct[4]), .B(ALUOp[1]), .C(n25), .D(n35), .Y(n18) );
  NOR2BX1 U5 ( .AN(ALUOp[1]), .B(n21), .Y(JumpR) );
  NAND2X1 U6 ( .A(n23), .B(n24), .Y(n26) );
  CLKINVX1 U7 ( .A(n25), .Y(n6) );
  CLKINVX1 U8 ( .A(n17), .Y(n8) );
  AND4X1 U9 ( .A(n7), .B(n35), .C(n10), .D(ALUOp[1]), .Y(Shift) );
  NOR3X1 U10 ( .A(n18), .B(funct[3]), .C(funct[1]), .Y(HI) );
  NOR3X1 U11 ( .A(n34), .B(funct[3]), .C(n18), .Y(LO) );
  OR2X1 U12 ( .A(JumpR), .B(raWrite), .Y(Jump) );
  NOR3X1 U13 ( .A(n34), .B(n7), .C(n18), .Y(Div) );
  NOR3X1 U14 ( .A(n18), .B(funct[1]), .C(n7), .Y(Mul) );
  NAND3BX1 U15 ( .AN(n11), .B(n12), .C(n13), .Y(RegWrite) );
  OAI31XL U16 ( .A0(n16), .A1(n6), .A2(n7), .B0(n8), .Y(n12) );
  NOR3BXL U17 ( .AN(n14), .B(inst[4]), .C(n15), .Y(n13) );
  NOR2X1 U18 ( .A(inst[4]), .B(n19), .Y(MemWrite) );
  NOR2BX1 U19 ( .AN(n22), .B(inst[4]), .Y(IF_Flush) );
  OAI222XL U20 ( .A0(n23), .A1(n5), .B0(eq), .B1(n24), .C0(n17), .C1(n21), .Y(
        n22) );
  CLKINVX1 U21 ( .A(eq), .Y(n5) );
  NOR2X1 U22 ( .A(n17), .B(inst[4]), .Y(ALUOp[1]) );
  NOR4X1 U23 ( .A(n32), .B(inst[1]), .C(inst[3]), .D(inst[5]), .Y(n29) );
  NOR2BX1 U24 ( .AN(n26), .B(inst[4]), .Y(Branch) );
  NAND4BX1 U25 ( .AN(inst[5]), .B(n9), .C(n32), .D(n27), .Y(n17) );
  NOR2X1 U26 ( .A(inst[1]), .B(inst[0]), .Y(n27) );
  NOR3X1 U27 ( .A(funct[1]), .B(funct[4]), .C(n6), .Y(n10) );
  NOR2X1 U28 ( .A(funct[5]), .B(funct[2]), .Y(n25) );
  NAND2BX1 U29 ( .AN(inst[0]), .B(n29), .Y(n23) );
  NAND2X1 U30 ( .A(n29), .B(inst[0]), .Y(n24) );
  NAND2X1 U31 ( .A(funct[3]), .B(n10), .Y(n21) );
  CLKINVX1 U32 ( .A(inst[3]), .Y(n9) );
  OAI221XL U33 ( .A0(n33), .A1(n32), .B0(inst[5]), .B1(n9), .C0(n30), .Y(n11)
         );
  AOI32X1 U34 ( .A0(n33), .A1(n32), .A2(inst[0]), .B0(inst[5]), .B1(n31), .Y(
        n30) );
  CLKINVX1 U35 ( .A(inst[1]), .Y(n33) );
  NOR2X1 U36 ( .A(n11), .B(n26), .Y(n28) );
  NOR3X1 U37 ( .A(inst[2]), .B(inst[3]), .C(n31), .Y(n20) );
  NOR2BX1 U38 ( .AN(n15), .B(inst[4]), .Y(raWrite) );
  NOR2BX1 U39 ( .AN(n20), .B(inst[5]), .Y(n15) );
  NAND4BX1 U40 ( .AN(n31), .B(inst[3]), .C(inst[5]), .D(n32), .Y(n19) );
  NAND2X1 U41 ( .A(inst[1]), .B(inst[0]), .Y(n31) );
  NAND2X1 U42 ( .A(inst[5]), .B(n20), .Y(n14) );
  CLKINVX1 U43 ( .A(funct[3]), .Y(n7) );
  CLKINVX1 U44 ( .A(funct[1]), .Y(n34) );
  CLKINVX1 U45 ( .A(funct[0]), .Y(n35) );
  NAND3BX1 U46 ( .AN(funct[4]), .B(n34), .C(n35), .Y(n16) );
  CLKBUFX3 U47 ( .A(IF_Flush), .Y(PCSrc) );
  CLKBUFX3 U48 ( .A(ALUOp[0]), .Y(ALURsc) );
  NAND4BX1 U49 ( .AN(inst[4]), .B(n19), .C(n14), .D(n28), .Y(ALUOp[0]) );
  CLKBUFX3 U50 ( .A(ALUOp[1]), .Y(RegDst) );
  CLKBUFX3 U51 ( .A(MemRead), .Y(MemtoReg) );
  NOR2X1 U52 ( .A(n14), .B(inst[4]), .Y(MemRead) );
endmodule


module BranchPrd ( clk, rst, taken, take, Branch );
  input clk, rst, taken, Branch;
  output take;
  wire   n2, n4, n5, n6, n7, n8, n1;
  wire   [1:0] state_r;

  DFFSX1 \state_r_reg[0]  ( .D(n8), .CK(clk), .SN(rst), .Q(state_r[0]), .QN(n2) );
  DFFSX1 \state_r_reg[1]  ( .D(n7), .CK(clk), .SN(rst), .Q(state_r[1]), .QN(
        take) );
  CLKINVX1 U3 ( .A(taken), .Y(n1) );
  OAI31XL U4 ( .A0(n4), .A1(taken), .A2(n2), .B0(n5), .Y(n7) );
  OAI31XL U5 ( .A0(n4), .A1(state_r[0]), .A2(n1), .B0(state_r[1]), .Y(n5) );
  NAND2X1 U6 ( .A(Branch), .B(n6), .Y(n4) );
  OAI222XL U7 ( .A0(state_r[1]), .A1(n2), .B0(taken), .B1(state_r[0]), .C0(
        take), .C1(n1), .Y(n6) );
  XOR2X1 U8 ( .A(n2), .B(n4), .Y(n8) );
endmodule


module forward_jump ( JumpR, Branch, RegJump, RegRt, IDEX_Opcode, 
        IDEX_RegWrite, IDEX_RegRt, IDEX_RegRd, EXMEM_RegWrite, EXMEM_MemRead, 
        EXMEM_RegRd, MEMWB_RegWrite, MEMWB_RegRd, ForwardJA, ForwardJB, stallJ
 );
  input [4:0] RegJump;
  input [4:0] RegRt;
  input [5:0] IDEX_Opcode;
  input [4:0] IDEX_RegRt;
  input [4:0] IDEX_RegRd;
  input [4:0] EXMEM_RegRd;
  input [4:0] MEMWB_RegRd;
  output [1:0] ForwardJA;
  output [1:0] ForwardJB;
  input JumpR, Branch, IDEX_RegWrite, EXMEM_RegWrite, EXMEM_MemRead,
         MEMWB_RegWrite;
  output stallJ;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;

  AOI2BB2X1 U2 ( .B0(n36), .B1(n37), .A0N(Branch), .A1N(JumpR), .Y(stallJ) );
  CLKINVX1 U3 ( .A(n88), .Y(ForwardJA[0]) );
  CLKINVX1 U4 ( .A(n75), .Y(ForwardJB[0]) );
  NOR4X1 U5 ( .A(n69), .B(n70), .C(n71), .D(n72), .Y(ForwardJB[1]) );
  XOR2X1 U6 ( .A(n3), .B(MEMWB_RegRd[2]), .Y(n70) );
  XOR2X1 U7 ( .A(n2), .B(MEMWB_RegRd[1]), .Y(n72) );
  XOR2X1 U8 ( .A(n1), .B(MEMWB_RegRd[0]), .Y(n71) );
  NOR4X1 U9 ( .A(n82), .B(n83), .C(n84), .D(n85), .Y(ForwardJA[1]) );
  XOR2X1 U10 ( .A(n8), .B(MEMWB_RegRd[2]), .Y(n83) );
  XOR2X1 U11 ( .A(n7), .B(MEMWB_RegRd[1]), .Y(n85) );
  XOR2X1 U12 ( .A(n6), .B(MEMWB_RegRd[0]), .Y(n84) );
  NOR2X1 U13 ( .A(n80), .B(n81), .Y(n78) );
  XOR2X1 U14 ( .A(n2), .B(EXMEM_RegRd[1]), .Y(n80) );
  XOR2X1 U15 ( .A(n5), .B(EXMEM_RegRd[4]), .Y(n81) );
  NAND4X1 U16 ( .A(n73), .B(n74), .C(MEMWB_RegWrite), .D(n75), .Y(n69) );
  XNOR2X1 U17 ( .A(MEMWB_RegRd[3]), .B(n4), .Y(n73) );
  XNOR2X1 U18 ( .A(MEMWB_RegRd[4]), .B(n5), .Y(n74) );
  NAND4X1 U19 ( .A(n86), .B(n87), .C(MEMWB_RegWrite), .D(n88), .Y(n82) );
  XNOR2X1 U20 ( .A(MEMWB_RegRd[3]), .B(n9), .Y(n86) );
  XNOR2X1 U21 ( .A(MEMWB_RegRd[4]), .B(n10), .Y(n87) );
  AND4X1 U22 ( .A(n89), .B(n90), .C(n91), .D(n92), .Y(n39) );
  XNOR2X1 U23 ( .A(EXMEM_RegRd[0]), .B(n6), .Y(n89) );
  XNOR2X1 U24 ( .A(EXMEM_RegRd[2]), .B(n8), .Y(n90) );
  XNOR2X1 U25 ( .A(EXMEM_RegRd[3]), .B(n9), .Y(n92) );
  AND4X1 U26 ( .A(n76), .B(n77), .C(n78), .D(n79), .Y(n38) );
  XNOR2X1 U27 ( .A(EXMEM_RegRd[0]), .B(n1), .Y(n76) );
  XNOR2X1 U28 ( .A(EXMEM_RegRd[2]), .B(n3), .Y(n77) );
  XNOR2X1 U29 ( .A(EXMEM_RegRd[3]), .B(n4), .Y(n79) );
  NAND3X1 U30 ( .A(n38), .B(n11), .C(EXMEM_RegWrite), .Y(n75) );
  NAND3X1 U31 ( .A(EXMEM_RegWrite), .B(n11), .C(n39), .Y(n88) );
  NOR2X1 U32 ( .A(n93), .B(n94), .Y(n91) );
  XOR2X1 U33 ( .A(n7), .B(EXMEM_RegRd[1]), .Y(n93) );
  XOR2X1 U34 ( .A(n10), .B(EXMEM_RegRd[4]), .Y(n94) );
  CLKBUFX3 U35 ( .A(RegRt[0]), .Y(n1) );
  CLKBUFX3 U36 ( .A(RegRt[2]), .Y(n3) );
  CLKBUFX3 U37 ( .A(RegJump[0]), .Y(n6) );
  CLKBUFX3 U38 ( .A(RegJump[2]), .Y(n8) );
  CLKBUFX3 U39 ( .A(RegRt[3]), .Y(n4) );
  CLKBUFX3 U40 ( .A(RegJump[3]), .Y(n9) );
  CLKBUFX3 U41 ( .A(RegRt[4]), .Y(n5) );
  CLKBUFX3 U42 ( .A(RegJump[4]), .Y(n10) );
  CLKBUFX3 U43 ( .A(RegRt[1]), .Y(n2) );
  CLKBUFX3 U44 ( .A(RegJump[1]), .Y(n7) );
  CLKINVX1 U45 ( .A(EXMEM_MemRead), .Y(n11) );
  NOR4X1 U46 ( .A(n49), .B(n50), .C(IDEX_Opcode[1]), .D(IDEX_Opcode[0]), .Y(
        n41) );
  OR4X1 U47 ( .A(IDEX_Opcode[3]), .B(IDEX_Opcode[2]), .C(IDEX_Opcode[5]), .D(
        IDEX_Opcode[4]), .Y(n49) );
  AOI33X1 U48 ( .A0(n51), .A1(n52), .A2(n53), .B0(n54), .B1(n55), .B2(n56), 
        .Y(n50) );
  XNOR2X1 U49 ( .A(IDEX_RegRd[0]), .B(n6), .Y(n51) );
  OAI21XL U50 ( .A0(n38), .A1(n39), .B0(EXMEM_MemRead), .Y(n37) );
  OAI31XL U51 ( .A0(n40), .A1(n41), .A2(n42), .B0(IDEX_RegWrite), .Y(n36) );
  NOR4X1 U52 ( .A(n63), .B(n64), .C(n65), .D(n66), .Y(n40) );
  XOR2X1 U53 ( .A(n5), .B(IDEX_RegRt[4]), .Y(n66) );
  XOR2X1 U54 ( .A(n2), .B(IDEX_RegRt[1]), .Y(n65) );
  XOR2X1 U55 ( .A(n4), .B(IDEX_RegRt[3]), .Y(n64) );
  XNOR2X1 U56 ( .A(IDEX_RegRd[2]), .B(n8), .Y(n52) );
  XNOR2X1 U57 ( .A(IDEX_RegRd[2]), .B(n3), .Y(n55) );
  XNOR2X1 U58 ( .A(IDEX_RegRd[0]), .B(n1), .Y(n54) );
  NOR4X1 U59 ( .A(n43), .B(n44), .C(n45), .D(n46), .Y(n42) );
  XOR2X1 U60 ( .A(n9), .B(IDEX_RegRt[3]), .Y(n44) );
  XOR2X1 U61 ( .A(n7), .B(IDEX_RegRt[1]), .Y(n45) );
  XOR2X1 U62 ( .A(n10), .B(IDEX_RegRt[4]), .Y(n46) );
  NOR3X1 U63 ( .A(n60), .B(n61), .C(n62), .Y(n53) );
  XOR2X1 U64 ( .A(n9), .B(IDEX_RegRd[3]), .Y(n60) );
  XOR2X1 U65 ( .A(n7), .B(IDEX_RegRd[1]), .Y(n61) );
  XOR2X1 U66 ( .A(n10), .B(IDEX_RegRd[4]), .Y(n62) );
  NOR3X1 U67 ( .A(n57), .B(n58), .C(n59), .Y(n56) );
  XOR2X1 U68 ( .A(n4), .B(IDEX_RegRd[3]), .Y(n57) );
  XOR2X1 U69 ( .A(n2), .B(IDEX_RegRd[1]), .Y(n58) );
  XOR2X1 U70 ( .A(n5), .B(IDEX_RegRd[4]), .Y(n59) );
  NAND2X1 U71 ( .A(n47), .B(n48), .Y(n43) );
  XNOR2X1 U72 ( .A(IDEX_RegRt[0]), .B(n6), .Y(n47) );
  XNOR2X1 U73 ( .A(IDEX_RegRt[2]), .B(n8), .Y(n48) );
  NAND2X1 U74 ( .A(n67), .B(n68), .Y(n63) );
  XNOR2X1 U75 ( .A(IDEX_RegRt[0]), .B(n1), .Y(n67) );
  XNOR2X1 U76 ( .A(IDEX_RegRt[2]), .B(n3), .Y(n68) );
endmodule


module HazardDetection ( opcode, IDEX_MemRead, IDEX_RegRt, IFID_RegRs, 
        IFID_RegRt, PCWrite, IFIDWrite, stall );
  input [5:0] opcode;
  input [4:0] IDEX_RegRt;
  input [4:0] IFID_RegRs;
  input [4:0] IFID_RegRt;
  input IDEX_MemRead;
  output PCWrite, IFIDWrite, stall;
  wire   n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29;

  OR4XL U3 ( .A(opcode[4]), .B(opcode[5]), .C(opcode[3]), .D(n29), .Y(n12) );
  NOR4XL U4 ( .A(n23), .B(opcode[3]), .C(opcode[5]), .D(opcode[4]), .Y(n20) );
  OAI31XL U5 ( .A0(n12), .A1(n13), .A2(n14), .B0(n15), .Y(stall) );
  NAND3X1 U6 ( .A(n27), .B(IDEX_MemRead), .C(n28), .Y(n13) );
  NAND3X1 U7 ( .A(n24), .B(n25), .C(n26), .Y(n14) );
  NAND4X1 U8 ( .A(n16), .B(n17), .C(n18), .D(n19), .Y(n15) );
  NOR4BX1 U9 ( .AN(IDEX_MemRead), .B(n20), .C(n21), .D(n22), .Y(n19) );
  XOR2X1 U10 ( .A(IFID_RegRs[4]), .B(IDEX_RegRt[4]), .Y(n21) );
  XOR2X1 U11 ( .A(IFID_RegRs[3]), .B(IDEX_RegRt[3]), .Y(n22) );
  XNOR2X1 U12 ( .A(IDEX_RegRt[2]), .B(IFID_RegRt[2]), .Y(n26) );
  XNOR2X1 U13 ( .A(IDEX_RegRt[4]), .B(IFID_RegRt[4]), .Y(n28) );
  XNOR2X1 U14 ( .A(IDEX_RegRt[0]), .B(IFID_RegRt[0]), .Y(n25) );
  XNOR2X1 U15 ( .A(IDEX_RegRt[1]), .B(IFID_RegRt[1]), .Y(n24) );
  XNOR2X1 U16 ( .A(IDEX_RegRt[3]), .B(IFID_RegRt[3]), .Y(n27) );
  NAND2BX1 U17 ( .AN(opcode[2]), .B(opcode[1]), .Y(n23) );
  OR3X2 U18 ( .A(opcode[0]), .B(opcode[2]), .C(opcode[1]), .Y(n29) );
  XNOR2X1 U19 ( .A(IDEX_RegRt[2]), .B(IFID_RegRs[2]), .Y(n18) );
  XNOR2X1 U20 ( .A(IDEX_RegRt[0]), .B(IFID_RegRs[0]), .Y(n17) );
  XNOR2X1 U21 ( .A(IDEX_RegRt[1]), .B(IFID_RegRs[1]), .Y(n16) );
  CLKBUFX3 U22 ( .A(PCWrite), .Y(IFIDWrite) );
  CLKINVX1 U23 ( .A(stall), .Y(PCWrite) );
endmodule


module register ( clk, rst_n, RegWrite, ReadReg1, ReadReg2, WriteReg, 
        WriteData, ReadData1, ReadData2 );
  input [4:0] ReadReg1;
  input [4:0] ReadReg2;
  input [4:0] WriteReg;
  input [31:0] WriteData;
  output [31:0] ReadData1;
  output [31:0] ReadData2;
  input clk, rst_n, RegWrite;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, \register_r[15][31] ,
         \register_r[15][30] , \register_r[15][29] , \register_r[15][28] ,
         \register_r[15][27] , \register_r[15][26] , \register_r[15][25] ,
         \register_r[15][24] , \register_r[15][23] , \register_r[15][22] ,
         \register_r[15][21] , \register_r[15][20] , \register_r[15][19] ,
         \register_r[15][18] , \register_r[15][17] , \register_r[15][16] ,
         \register_r[15][15] , \register_r[15][14] , \register_r[15][13] ,
         \register_r[15][12] , \register_r[15][11] , \register_r[15][10] ,
         \register_r[15][9] , \register_r[15][8] , \register_r[15][7] ,
         \register_r[15][6] , \register_r[15][5] , \register_r[15][4] ,
         \register_r[15][3] , \register_r[15][2] , \register_r[15][1] ,
         \register_r[15][0] , \register_r[14][31] , \register_r[14][30] ,
         \register_r[14][29] , \register_r[14][28] , \register_r[14][27] ,
         \register_r[14][26] , \register_r[14][25] , \register_r[14][24] ,
         \register_r[14][23] , \register_r[14][22] , \register_r[14][21] ,
         \register_r[14][20] , \register_r[14][19] , \register_r[14][18] ,
         \register_r[14][17] , \register_r[14][16] , \register_r[14][15] ,
         \register_r[14][14] , \register_r[14][13] , \register_r[14][12] ,
         \register_r[14][11] , \register_r[14][10] , \register_r[14][9] ,
         \register_r[14][8] , \register_r[14][7] , \register_r[14][6] ,
         \register_r[14][5] , \register_r[14][4] , \register_r[14][3] ,
         \register_r[14][2] , \register_r[14][1] , \register_r[14][0] ,
         \register_r[11][31] , \register_r[11][30] , \register_r[11][29] ,
         \register_r[11][28] , \register_r[11][27] , \register_r[11][26] ,
         \register_r[11][25] , \register_r[11][24] , \register_r[11][23] ,
         \register_r[11][22] , \register_r[11][21] , \register_r[11][20] ,
         \register_r[11][19] , \register_r[11][18] , \register_r[11][17] ,
         \register_r[11][16] , \register_r[11][15] , \register_r[11][14] ,
         \register_r[11][13] , \register_r[11][12] , \register_r[11][11] ,
         \register_r[11][10] , \register_r[11][9] , \register_r[11][8] ,
         \register_r[11][7] , \register_r[11][6] , \register_r[11][5] ,
         \register_r[11][4] , \register_r[11][3] , \register_r[11][2] ,
         \register_r[11][1] , \register_r[11][0] , \register_r[10][31] ,
         \register_r[10][30] , \register_r[10][29] , \register_r[10][28] ,
         \register_r[10][27] , \register_r[10][26] , \register_r[10][25] ,
         \register_r[10][24] , \register_r[10][23] , \register_r[10][22] ,
         \register_r[10][21] , \register_r[10][20] , \register_r[10][19] ,
         \register_r[10][18] , \register_r[10][17] , \register_r[10][16] ,
         \register_r[10][15] , \register_r[10][14] , \register_r[10][13] ,
         \register_r[10][12] , \register_r[10][11] , \register_r[10][10] ,
         \register_r[10][9] , \register_r[10][8] , \register_r[10][7] ,
         \register_r[10][6] , \register_r[10][5] , \register_r[10][4] ,
         \register_r[10][3] , \register_r[10][2] , \register_r[10][1] ,
         \register_r[10][0] , \register_r[9][31] , \register_r[9][30] ,
         \register_r[9][29] , \register_r[9][28] , \register_r[9][27] ,
         \register_r[9][26] , \register_r[9][25] , \register_r[9][24] ,
         \register_r[9][23] , \register_r[9][22] , \register_r[9][21] ,
         \register_r[9][20] , \register_r[9][19] , \register_r[9][18] ,
         \register_r[9][17] , \register_r[9][16] , \register_r[9][15] ,
         \register_r[9][14] , \register_r[9][13] , \register_r[9][12] ,
         \register_r[9][11] , \register_r[9][10] , \register_r[9][9] ,
         \register_r[9][8] , \register_r[9][7] , \register_r[9][6] ,
         \register_r[9][5] , \register_r[9][4] , \register_r[9][3] ,
         \register_r[9][2] , \register_r[9][1] , \register_r[9][0] ,
         \register_r[8][31] , \register_r[8][30] , \register_r[8][29] ,
         \register_r[8][28] , \register_r[8][27] , \register_r[8][26] ,
         \register_r[8][25] , \register_r[8][24] , \register_r[8][23] ,
         \register_r[8][22] , \register_r[8][21] , \register_r[8][20] ,
         \register_r[8][19] , \register_r[8][18] , \register_r[8][17] ,
         \register_r[8][16] , \register_r[8][15] , \register_r[8][14] ,
         \register_r[8][13] , \register_r[8][12] , \register_r[8][11] ,
         \register_r[8][10] , \register_r[8][9] , \register_r[8][8] ,
         \register_r[8][7] , \register_r[8][6] , \register_r[8][5] ,
         \register_r[8][4] , \register_r[8][3] , \register_r[8][2] ,
         \register_r[8][1] , \register_r[8][0] , \register_r[7][31] ,
         \register_r[7][30] , \register_r[7][29] , \register_r[7][28] ,
         \register_r[7][27] , \register_r[7][26] , \register_r[7][25] ,
         \register_r[7][24] , \register_r[7][23] , \register_r[7][22] ,
         \register_r[7][21] , \register_r[7][20] , \register_r[7][19] ,
         \register_r[7][18] , \register_r[7][17] , \register_r[7][16] ,
         \register_r[7][15] , \register_r[7][14] , \register_r[7][13] ,
         \register_r[7][12] , \register_r[7][11] , \register_r[7][10] ,
         \register_r[7][9] , \register_r[7][8] , \register_r[7][7] ,
         \register_r[7][6] , \register_r[7][5] , \register_r[7][4] ,
         \register_r[7][3] , \register_r[7][2] , \register_r[7][1] ,
         \register_r[7][0] , \register_r[6][31] , \register_r[6][30] ,
         \register_r[6][29] , \register_r[6][28] , \register_r[6][27] ,
         \register_r[6][26] , \register_r[6][25] , \register_r[6][24] ,
         \register_r[6][23] , \register_r[6][22] , \register_r[6][21] ,
         \register_r[6][20] , \register_r[6][19] , \register_r[6][18] ,
         \register_r[6][17] , \register_r[6][16] , \register_r[6][15] ,
         \register_r[6][14] , \register_r[6][13] , \register_r[6][12] ,
         \register_r[6][11] , \register_r[6][10] , \register_r[6][9] ,
         \register_r[6][8] , \register_r[6][7] , \register_r[6][6] ,
         \register_r[6][5] , \register_r[6][4] , \register_r[6][3] ,
         \register_r[6][2] , \register_r[6][1] , \register_r[6][0] ,
         \register_r[5][31] , \register_r[5][30] , \register_r[5][29] ,
         \register_r[5][28] , \register_r[5][27] , \register_r[5][26] ,
         \register_r[5][25] , \register_r[5][24] , \register_r[5][23] ,
         \register_r[5][22] , \register_r[5][21] , \register_r[5][20] ,
         \register_r[5][19] , \register_r[5][18] , \register_r[5][17] ,
         \register_r[5][16] , \register_r[5][15] , \register_r[5][14] ,
         \register_r[5][13] , \register_r[5][12] , \register_r[5][11] ,
         \register_r[5][10] , \register_r[5][9] , \register_r[5][8] ,
         \register_r[5][7] , \register_r[5][6] , \register_r[5][5] ,
         \register_r[5][4] , \register_r[5][3] , \register_r[5][2] ,
         \register_r[5][1] , \register_r[5][0] , \register_r[4][31] ,
         \register_r[4][30] , \register_r[4][29] , \register_r[4][28] ,
         \register_r[4][27] , \register_r[4][26] , \register_r[4][25] ,
         \register_r[4][24] , \register_r[4][23] , \register_r[4][22] ,
         \register_r[4][21] , \register_r[4][20] , \register_r[4][19] ,
         \register_r[4][18] , \register_r[4][17] , \register_r[4][16] ,
         \register_r[4][15] , \register_r[4][14] , \register_r[4][13] ,
         \register_r[4][12] , \register_r[4][11] , \register_r[4][10] ,
         \register_r[4][9] , \register_r[4][8] , \register_r[4][7] ,
         \register_r[4][6] , \register_r[4][5] , \register_r[4][4] ,
         \register_r[4][3] , \register_r[4][2] , \register_r[4][1] ,
         \register_r[4][0] , \register_r[3][31] , \register_r[3][30] ,
         \register_r[3][29] , \register_r[3][28] , \register_r[3][27] ,
         \register_r[3][26] , \register_r[3][25] , \register_r[3][24] ,
         \register_r[3][23] , \register_r[3][22] , \register_r[3][21] ,
         \register_r[3][20] , \register_r[3][19] , \register_r[3][18] ,
         \register_r[3][17] , \register_r[3][16] , \register_r[3][15] ,
         \register_r[3][14] , \register_r[3][13] , \register_r[3][12] ,
         \register_r[3][11] , \register_r[3][10] , \register_r[3][9] ,
         \register_r[3][8] , \register_r[3][7] , \register_r[3][6] ,
         \register_r[3][5] , \register_r[3][4] , \register_r[3][3] ,
         \register_r[3][2] , \register_r[3][1] , \register_r[3][0] ,
         \register_r[1][31] , \register_r[1][30] , \register_r[1][29] ,
         \register_r[1][28] , \register_r[1][27] , \register_r[1][26] ,
         \register_r[1][25] , \register_r[1][24] , \register_r[1][23] ,
         \register_r[1][22] , \register_r[1][21] , \register_r[1][20] ,
         \register_r[1][19] , \register_r[1][18] , \register_r[1][17] ,
         \register_r[1][16] , \register_r[1][15] , \register_r[1][14] ,
         \register_r[1][13] , \register_r[1][12] , \register_r[1][11] ,
         \register_r[1][10] , \register_r[1][9] , \register_r[1][8] ,
         \register_r[1][7] , \register_r[1][6] , \register_r[1][5] ,
         \register_r[1][4] , \register_r[1][3] , \register_r[1][2] ,
         \register_r[1][1] , \register_r[1][0] , \register_r[31][31] ,
         \register_r[31][30] , \register_r[31][29] , \register_r[31][28] ,
         \register_r[31][27] , \register_r[31][26] , \register_r[31][25] ,
         \register_r[31][24] , \register_r[31][23] , \register_r[31][22] ,
         \register_r[31][21] , \register_r[31][20] , \register_r[31][19] ,
         \register_r[31][18] , \register_r[31][17] , \register_r[31][16] ,
         \register_r[31][15] , \register_r[31][14] , \register_r[31][13] ,
         \register_r[31][12] , \register_r[31][11] , \register_r[31][10] ,
         \register_r[31][9] , \register_r[31][8] , \register_r[31][7] ,
         \register_r[31][6] , \register_r[31][5] , \register_r[31][4] ,
         \register_r[31][3] , \register_r[31][2] , \register_r[31][1] ,
         \register_r[31][0] , \register_r[30][31] , \register_r[30][30] ,
         \register_r[30][29] , \register_r[30][28] , \register_r[30][27] ,
         \register_r[30][26] , \register_r[30][25] , \register_r[30][24] ,
         \register_r[30][23] , \register_r[30][22] , \register_r[30][21] ,
         \register_r[30][20] , \register_r[30][19] , \register_r[30][18] ,
         \register_r[30][17] , \register_r[30][16] , \register_r[30][15] ,
         \register_r[30][14] , \register_r[30][13] , \register_r[30][12] ,
         \register_r[30][11] , \register_r[30][10] , \register_r[30][9] ,
         \register_r[30][8] , \register_r[30][7] , \register_r[30][6] ,
         \register_r[30][5] , \register_r[30][4] , \register_r[30][3] ,
         \register_r[30][2] , \register_r[30][1] , \register_r[30][0] ,
         \register_r[29][31] , \register_r[29][30] , \register_r[29][29] ,
         \register_r[29][28] , \register_r[29][27] , \register_r[29][26] ,
         \register_r[29][25] , \register_r[29][24] , \register_r[29][23] ,
         \register_r[29][22] , \register_r[29][21] , \register_r[29][20] ,
         \register_r[29][19] , \register_r[29][18] , \register_r[29][17] ,
         \register_r[29][16] , \register_r[29][15] , \register_r[29][14] ,
         \register_r[29][13] , \register_r[29][12] , \register_r[29][11] ,
         \register_r[29][10] , \register_r[29][9] , \register_r[29][8] ,
         \register_r[29][7] , \register_r[29][6] , \register_r[29][5] ,
         \register_r[29][4] , \register_r[29][3] , \register_r[29][2] ,
         \register_r[29][1] , \register_r[29][0] , \register_r[28][31] ,
         \register_r[28][30] , \register_r[28][29] , \register_r[28][28] ,
         \register_r[28][27] , \register_r[28][26] , \register_r[28][25] ,
         \register_r[28][24] , \register_r[28][23] , \register_r[28][22] ,
         \register_r[28][21] , \register_r[28][20] , \register_r[28][19] ,
         \register_r[28][18] , \register_r[28][17] , \register_r[28][16] ,
         \register_r[28][15] , \register_r[28][14] , \register_r[28][13] ,
         \register_r[28][12] , \register_r[28][11] , \register_r[28][10] ,
         \register_r[28][9] , \register_r[28][8] , \register_r[28][7] ,
         \register_r[28][6] , \register_r[28][5] , \register_r[28][4] ,
         \register_r[28][3] , \register_r[28][2] , \register_r[28][1] ,
         \register_r[28][0] , \register_r[27][31] , \register_r[27][30] ,
         \register_r[27][29] , \register_r[27][28] , \register_r[27][27] ,
         \register_r[27][26] , \register_r[27][25] , \register_r[27][24] ,
         \register_r[27][23] , \register_r[27][22] , \register_r[27][21] ,
         \register_r[27][20] , \register_r[27][19] , \register_r[27][18] ,
         \register_r[27][17] , \register_r[27][16] , \register_r[27][15] ,
         \register_r[27][14] , \register_r[27][13] , \register_r[27][12] ,
         \register_r[27][11] , \register_r[27][10] , \register_r[27][9] ,
         \register_r[27][8] , \register_r[27][7] , \register_r[27][6] ,
         \register_r[27][5] , \register_r[27][4] , \register_r[27][3] ,
         \register_r[27][2] , \register_r[27][1] , \register_r[27][0] ,
         \register_r[26][31] , \register_r[26][30] , \register_r[26][29] ,
         \register_r[26][28] , \register_r[26][27] , \register_r[26][26] ,
         \register_r[26][25] , \register_r[26][24] , \register_r[26][23] ,
         \register_r[26][22] , \register_r[26][21] , \register_r[26][20] ,
         \register_r[26][19] , \register_r[26][18] , \register_r[26][17] ,
         \register_r[26][16] , \register_r[26][15] , \register_r[26][14] ,
         \register_r[26][13] , \register_r[26][12] , \register_r[26][11] ,
         \register_r[26][10] , \register_r[26][9] , \register_r[26][8] ,
         \register_r[26][7] , \register_r[26][6] , \register_r[26][5] ,
         \register_r[26][4] , \register_r[26][3] , \register_r[26][2] ,
         \register_r[26][1] , \register_r[26][0] , \register_r[25][31] ,
         \register_r[25][30] , \register_r[25][29] , \register_r[25][28] ,
         \register_r[25][27] , \register_r[25][26] , \register_r[25][25] ,
         \register_r[25][24] , \register_r[25][23] , \register_r[25][22] ,
         \register_r[25][21] , \register_r[25][20] , \register_r[25][19] ,
         \register_r[25][18] , \register_r[25][17] , \register_r[25][16] ,
         \register_r[25][15] , \register_r[25][14] , \register_r[25][13] ,
         \register_r[25][12] , \register_r[25][11] , \register_r[25][10] ,
         \register_r[25][9] , \register_r[25][8] , \register_r[25][7] ,
         \register_r[25][6] , \register_r[25][5] , \register_r[25][4] ,
         \register_r[25][3] , \register_r[25][2] , \register_r[25][1] ,
         \register_r[25][0] , \register_r[24][31] , \register_r[24][30] ,
         \register_r[24][29] , \register_r[24][28] , \register_r[24][27] ,
         \register_r[24][26] , \register_r[24][25] , \register_r[24][24] ,
         \register_r[24][23] , \register_r[24][22] , \register_r[24][21] ,
         \register_r[24][20] , \register_r[24][19] , \register_r[24][18] ,
         \register_r[24][17] , \register_r[24][16] , \register_r[24][15] ,
         \register_r[24][14] , \register_r[24][13] , \register_r[24][12] ,
         \register_r[24][11] , \register_r[24][10] , \register_r[24][9] ,
         \register_r[24][8] , \register_r[24][7] , \register_r[24][6] ,
         \register_r[24][5] , \register_r[24][4] , \register_r[24][3] ,
         \register_r[24][2] , \register_r[24][1] , \register_r[24][0] ,
         \register_r[23][31] , \register_r[23][30] , \register_r[23][29] ,
         \register_r[23][28] , \register_r[23][27] , \register_r[23][26] ,
         \register_r[23][25] , \register_r[23][24] , \register_r[23][23] ,
         \register_r[23][22] , \register_r[23][21] , \register_r[23][20] ,
         \register_r[23][19] , \register_r[23][18] , \register_r[23][17] ,
         \register_r[23][16] , \register_r[23][15] , \register_r[23][14] ,
         \register_r[23][13] , \register_r[23][12] , \register_r[23][11] ,
         \register_r[23][10] , \register_r[23][9] , \register_r[23][8] ,
         \register_r[23][7] , \register_r[23][6] , \register_r[23][5] ,
         \register_r[23][4] , \register_r[23][3] , \register_r[23][2] ,
         \register_r[23][1] , \register_r[23][0] , \register_r[22][31] ,
         \register_r[22][30] , \register_r[22][29] , \register_r[22][28] ,
         \register_r[22][27] , \register_r[22][26] , \register_r[22][25] ,
         \register_r[22][24] , \register_r[22][23] , \register_r[22][22] ,
         \register_r[22][21] , \register_r[22][20] , \register_r[22][19] ,
         \register_r[22][18] , \register_r[22][17] , \register_r[22][16] ,
         \register_r[22][15] , \register_r[22][14] , \register_r[22][13] ,
         \register_r[22][12] , \register_r[22][11] , \register_r[22][10] ,
         \register_r[22][9] , \register_r[22][8] , \register_r[22][7] ,
         \register_r[22][6] , \register_r[22][5] , \register_r[22][4] ,
         \register_r[22][3] , \register_r[22][2] , \register_r[22][1] ,
         \register_r[22][0] , \register_r[21][31] , \register_r[21][30] ,
         \register_r[21][29] , \register_r[21][28] , \register_r[21][27] ,
         \register_r[21][26] , \register_r[21][25] , \register_r[21][24] ,
         \register_r[21][23] , \register_r[21][22] , \register_r[21][21] ,
         \register_r[21][20] , \register_r[21][19] , \register_r[21][18] ,
         \register_r[21][17] , \register_r[21][16] , \register_r[21][15] ,
         \register_r[21][14] , \register_r[21][13] , \register_r[21][12] ,
         \register_r[21][11] , \register_r[21][10] , \register_r[21][9] ,
         \register_r[21][8] , \register_r[21][7] , \register_r[21][6] ,
         \register_r[21][5] , \register_r[21][4] , \register_r[21][3] ,
         \register_r[21][2] , \register_r[21][1] , \register_r[21][0] ,
         \register_r[20][31] , \register_r[20][30] , \register_r[20][29] ,
         \register_r[20][28] , \register_r[20][27] , \register_r[20][26] ,
         \register_r[20][25] , \register_r[20][24] , \register_r[20][23] ,
         \register_r[20][22] , \register_r[20][21] , \register_r[20][20] ,
         \register_r[20][19] , \register_r[20][18] , \register_r[20][17] ,
         \register_r[20][16] , \register_r[20][15] , \register_r[20][14] ,
         \register_r[20][13] , \register_r[20][12] , \register_r[20][11] ,
         \register_r[20][10] , \register_r[20][9] , \register_r[20][8] ,
         \register_r[20][7] , \register_r[20][6] , \register_r[20][5] ,
         \register_r[20][4] , \register_r[20][3] , \register_r[20][2] ,
         \register_r[20][1] , \register_r[20][0] , \register_r[19][31] ,
         \register_r[19][30] , \register_r[19][29] , \register_r[19][28] ,
         \register_r[19][27] , \register_r[19][26] , \register_r[19][25] ,
         \register_r[19][24] , \register_r[19][23] , \register_r[19][22] ,
         \register_r[19][21] , \register_r[19][20] , \register_r[19][19] ,
         \register_r[19][18] , \register_r[19][17] , \register_r[19][16] ,
         \register_r[19][15] , \register_r[19][14] , \register_r[19][13] ,
         \register_r[19][12] , \register_r[19][11] , \register_r[19][10] ,
         \register_r[19][9] , \register_r[19][8] , \register_r[19][7] ,
         \register_r[19][6] , \register_r[19][5] , \register_r[19][4] ,
         \register_r[19][3] , \register_r[19][2] , \register_r[19][1] ,
         \register_r[19][0] , \register_r[18][31] , \register_r[18][30] ,
         \register_r[18][29] , \register_r[18][28] , \register_r[18][27] ,
         \register_r[18][26] , \register_r[18][25] , \register_r[18][24] ,
         \register_r[18][23] , \register_r[18][22] , \register_r[18][21] ,
         \register_r[18][20] , \register_r[18][19] , \register_r[18][18] ,
         \register_r[18][17] , \register_r[18][16] , \register_r[18][15] ,
         \register_r[18][14] , \register_r[18][13] , \register_r[18][12] ,
         \register_r[18][11] , \register_r[18][10] , \register_r[18][9] ,
         \register_r[18][8] , \register_r[18][7] , \register_r[18][6] ,
         \register_r[18][5] , \register_r[18][4] , \register_r[18][3] ,
         \register_r[18][2] , \register_r[18][1] , \register_r[18][0] ,
         \register_r[17][31] , \register_r[17][30] , \register_r[17][29] ,
         \register_r[17][28] , \register_r[17][27] , \register_r[17][26] ,
         \register_r[17][25] , \register_r[17][24] , \register_r[17][23] ,
         \register_r[17][22] , \register_r[17][21] , \register_r[17][20] ,
         \register_r[17][19] , \register_r[17][18] , \register_r[17][17] ,
         \register_r[17][16] , \register_r[17][15] , \register_r[17][14] ,
         \register_r[17][13] , \register_r[17][12] , \register_r[17][11] ,
         \register_r[17][10] , \register_r[17][9] , \register_r[17][8] ,
         \register_r[17][7] , \register_r[17][6] , \register_r[17][5] ,
         \register_r[17][4] , \register_r[17][3] , \register_r[17][2] ,
         \register_r[17][1] , \register_r[17][0] , \register_r[16][31] ,
         \register_r[16][30] , \register_r[16][29] , \register_r[16][28] ,
         \register_r[16][27] , \register_r[16][26] , \register_r[16][25] ,
         \register_r[16][24] , \register_r[16][23] , \register_r[16][22] ,
         \register_r[16][21] , \register_r[16][20] , \register_r[16][19] ,
         \register_r[16][18] , \register_r[16][17] , \register_r[16][16] ,
         \register_r[16][15] , \register_r[16][14] , \register_r[16][13] ,
         \register_r[16][12] , \register_r[16][11] , \register_r[16][10] ,
         \register_r[16][9] , \register_r[16][8] , \register_r[16][7] ,
         \register_r[16][6] , \register_r[16][5] , \register_r[16][4] ,
         \register_r[16][3] , \register_r[16][2] , \register_r[16][1] ,
         \register_r[16][0] , n9, n43, n44, n45, n47, n48, n49, n51, n53, n54,
         n56, n58, n59, n60, n64, n66, n67, n69, n70, n72, n74, n76, n78, n80,
         n81, n84, n86, n87, n89, n90, n92, n94, n96, n98, n100, n101, n103,
         n104, n106, n107, n109, n110, n112, n115, n117, n120, n122, n123,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n1, n2, n3,
         n4, n5, n6, n7, n8, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n46, n50, n52, n55, n57,
         n61, n62, n63, n65, n68, n71, n73, n75, n77, n79, n82, n83, n85, n88,
         n91, n93, n95, n97, n99, n102, n105, n108, n111, n113, n114, n116,
         n118, n119, n121, n124, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444;
  wire   [31:0] r_12;
  wire   [31:0] r_13;
  wire   [31:0] prev_ReadData1;
  wire   [31:0] prev_ReadData2;
  assign N2 = ReadReg1[0];
  assign N3 = ReadReg1[1];
  assign N4 = ReadReg1[2];
  assign N5 = ReadReg1[3];
  assign N6 = ReadReg1[4];
  assign N7 = ReadReg2[0];
  assign N8 = ReadReg2[1];
  assign N9 = ReadReg2[2];
  assign N10 = ReadReg2[3];
  assign N11 = ReadReg2[4];

  DFFRX1 \register_r_reg[31][31]  ( .D(n2122), .CK(clk), .RN(n3381), .Q(
        \register_r[31][31] ), .QN(n139) );
  DFFRX1 \register_r_reg[31][30]  ( .D(n2121), .CK(clk), .RN(n3381), .Q(
        \register_r[31][30] ), .QN(n140) );
  DFFRX1 \register_r_reg[31][29]  ( .D(n2120), .CK(clk), .RN(n3381), .Q(
        \register_r[31][29] ), .QN(n141) );
  DFFRX1 \register_r_reg[31][28]  ( .D(n2119), .CK(clk), .RN(n3381), .Q(
        \register_r[31][28] ), .QN(n142) );
  DFFRX1 \register_r_reg[31][27]  ( .D(n2118), .CK(clk), .RN(n3381), .Q(
        \register_r[31][27] ), .QN(n143) );
  DFFRX1 \register_r_reg[31][26]  ( .D(n2117), .CK(clk), .RN(n3381), .Q(
        \register_r[31][26] ), .QN(n144) );
  DFFRX1 \register_r_reg[31][25]  ( .D(n2116), .CK(clk), .RN(n3381), .Q(
        \register_r[31][25] ), .QN(n145) );
  DFFRX1 \register_r_reg[31][24]  ( .D(n2115), .CK(clk), .RN(n3381), .Q(
        \register_r[31][24] ), .QN(n146) );
  DFFRX1 \register_r_reg[31][23]  ( .D(n2114), .CK(clk), .RN(n3380), .Q(
        \register_r[31][23] ), .QN(n147) );
  DFFRX1 \register_r_reg[31][22]  ( .D(n2113), .CK(clk), .RN(n3380), .Q(
        \register_r[31][22] ), .QN(n148) );
  DFFRX1 \register_r_reg[31][21]  ( .D(n2112), .CK(clk), .RN(n3380), .Q(
        \register_r[31][21] ), .QN(n149) );
  DFFRX1 \register_r_reg[31][20]  ( .D(n2111), .CK(clk), .RN(n3380), .Q(
        \register_r[31][20] ), .QN(n150) );
  DFFRX1 \register_r_reg[31][19]  ( .D(n2110), .CK(clk), .RN(n3380), .Q(
        \register_r[31][19] ), .QN(n151) );
  DFFRX1 \register_r_reg[31][18]  ( .D(n2109), .CK(clk), .RN(n3380), .Q(
        \register_r[31][18] ), .QN(n152) );
  DFFRX1 \register_r_reg[31][17]  ( .D(n2108), .CK(clk), .RN(n3380), .Q(
        \register_r[31][17] ), .QN(n153) );
  DFFRX1 \register_r_reg[31][16]  ( .D(n2107), .CK(clk), .RN(n3380), .Q(
        \register_r[31][16] ), .QN(n154) );
  DFFRX1 \register_r_reg[31][15]  ( .D(n2106), .CK(clk), .RN(n3380), .Q(
        \register_r[31][15] ), .QN(n155) );
  DFFRX1 \register_r_reg[31][14]  ( .D(n2105), .CK(clk), .RN(n3380), .Q(
        \register_r[31][14] ), .QN(n156) );
  DFFRX1 \register_r_reg[31][13]  ( .D(n2104), .CK(clk), .RN(n3380), .Q(
        \register_r[31][13] ), .QN(n157) );
  DFFRX1 \register_r_reg[31][12]  ( .D(n2103), .CK(clk), .RN(n3380), .Q(
        \register_r[31][12] ), .QN(n158) );
  DFFRX1 \register_r_reg[31][11]  ( .D(n2102), .CK(clk), .RN(n3379), .Q(
        \register_r[31][11] ), .QN(n159) );
  DFFRX1 \register_r_reg[31][10]  ( .D(n2101), .CK(clk), .RN(n3379), .Q(
        \register_r[31][10] ), .QN(n160) );
  DFFRX1 \register_r_reg[31][9]  ( .D(n2100), .CK(clk), .RN(n3379), .Q(
        \register_r[31][9] ), .QN(n161) );
  DFFRX1 \register_r_reg[31][8]  ( .D(n2099), .CK(clk), .RN(n3379), .Q(
        \register_r[31][8] ), .QN(n162) );
  DFFRX1 \register_r_reg[31][7]  ( .D(n2098), .CK(clk), .RN(n3379), .Q(
        \register_r[31][7] ), .QN(n163) );
  DFFRX1 \register_r_reg[31][6]  ( .D(n2097), .CK(clk), .RN(n3379), .Q(
        \register_r[31][6] ), .QN(n164) );
  DFFRX1 \register_r_reg[31][5]  ( .D(n2096), .CK(clk), .RN(n3379), .Q(
        \register_r[31][5] ), .QN(n165) );
  DFFRX1 \register_r_reg[31][4]  ( .D(n2095), .CK(clk), .RN(n3379), .Q(
        \register_r[31][4] ), .QN(n166) );
  DFFRX1 \register_r_reg[31][3]  ( .D(n2094), .CK(clk), .RN(n3379), .Q(
        \register_r[31][3] ), .QN(n167) );
  DFFRX1 \register_r_reg[31][2]  ( .D(n2093), .CK(clk), .RN(n3379), .Q(
        \register_r[31][2] ), .QN(n168) );
  DFFRX1 \register_r_reg[31][1]  ( .D(n2092), .CK(clk), .RN(n3379), .Q(
        \register_r[31][1] ), .QN(n169) );
  DFFRX1 \register_r_reg[31][0]  ( .D(n2091), .CK(clk), .RN(n3379), .Q(
        \register_r[31][0] ), .QN(n170) );
  DFFRX1 \register_r_reg[27][31]  ( .D(n1994), .CK(clk), .RN(n3370), .Q(
        \register_r[27][31] ), .QN(n267) );
  DFFRX1 \register_r_reg[27][30]  ( .D(n1993), .CK(clk), .RN(n3370), .Q(
        \register_r[27][30] ), .QN(n268) );
  DFFRX1 \register_r_reg[27][29]  ( .D(n1992), .CK(clk), .RN(n3370), .Q(
        \register_r[27][29] ), .QN(n269) );
  DFFRX1 \register_r_reg[27][28]  ( .D(n1991), .CK(clk), .RN(n3370), .Q(
        \register_r[27][28] ), .QN(n270) );
  DFFRX1 \register_r_reg[27][27]  ( .D(n1990), .CK(clk), .RN(n3370), .Q(
        \register_r[27][27] ), .QN(n271) );
  DFFRX1 \register_r_reg[27][26]  ( .D(n1989), .CK(clk), .RN(n3370), .Q(
        \register_r[27][26] ), .QN(n272) );
  DFFRX1 \register_r_reg[27][25]  ( .D(n1988), .CK(clk), .RN(n3370), .Q(
        \register_r[27][25] ), .QN(n273) );
  DFFRX1 \register_r_reg[27][24]  ( .D(n1987), .CK(clk), .RN(n3370), .Q(
        \register_r[27][24] ), .QN(n274) );
  DFFRX1 \register_r_reg[27][23]  ( .D(n1986), .CK(clk), .RN(n3370), .Q(
        \register_r[27][23] ), .QN(n275) );
  DFFRX1 \register_r_reg[27][22]  ( .D(n1985), .CK(clk), .RN(n3370), .Q(
        \register_r[27][22] ), .QN(n276) );
  DFFRX1 \register_r_reg[27][21]  ( .D(n1984), .CK(clk), .RN(n3370), .Q(
        \register_r[27][21] ), .QN(n277) );
  DFFRX1 \register_r_reg[27][20]  ( .D(n1983), .CK(clk), .RN(n3370), .Q(
        \register_r[27][20] ), .QN(n278) );
  DFFRX1 \register_r_reg[27][19]  ( .D(n1982), .CK(clk), .RN(n3369), .Q(
        \register_r[27][19] ), .QN(n279) );
  DFFRX1 \register_r_reg[27][18]  ( .D(n1981), .CK(clk), .RN(n3369), .Q(
        \register_r[27][18] ), .QN(n280) );
  DFFRX1 \register_r_reg[27][17]  ( .D(n1980), .CK(clk), .RN(n3369), .Q(
        \register_r[27][17] ), .QN(n281) );
  DFFRX1 \register_r_reg[27][16]  ( .D(n1979), .CK(clk), .RN(n3369), .Q(
        \register_r[27][16] ), .QN(n282) );
  DFFRX1 \register_r_reg[27][15]  ( .D(n1978), .CK(clk), .RN(n3369), .Q(
        \register_r[27][15] ), .QN(n283) );
  DFFRX1 \register_r_reg[27][14]  ( .D(n1977), .CK(clk), .RN(n3369), .Q(
        \register_r[27][14] ), .QN(n284) );
  DFFRX1 \register_r_reg[27][13]  ( .D(n1976), .CK(clk), .RN(n3369), .Q(
        \register_r[27][13] ), .QN(n285) );
  DFFRX1 \register_r_reg[27][12]  ( .D(n1975), .CK(clk), .RN(n3369), .Q(
        \register_r[27][12] ), .QN(n286) );
  DFFRX1 \register_r_reg[27][11]  ( .D(n1974), .CK(clk), .RN(n3369), .Q(
        \register_r[27][11] ), .QN(n287) );
  DFFRX1 \register_r_reg[27][10]  ( .D(n1973), .CK(clk), .RN(n3369), .Q(
        \register_r[27][10] ), .QN(n288) );
  DFFRX1 \register_r_reg[27][9]  ( .D(n1972), .CK(clk), .RN(n3369), .Q(
        \register_r[27][9] ), .QN(n289) );
  DFFRX1 \register_r_reg[27][8]  ( .D(n1971), .CK(clk), .RN(n3369), .Q(
        \register_r[27][8] ), .QN(n290) );
  DFFRX1 \register_r_reg[27][7]  ( .D(n1970), .CK(clk), .RN(n3368), .Q(
        \register_r[27][7] ), .QN(n291) );
  DFFRX1 \register_r_reg[27][6]  ( .D(n1969), .CK(clk), .RN(n3368), .Q(
        \register_r[27][6] ), .QN(n292) );
  DFFRX1 \register_r_reg[27][5]  ( .D(n1968), .CK(clk), .RN(n3368), .Q(
        \register_r[27][5] ), .QN(n293) );
  DFFRX1 \register_r_reg[27][4]  ( .D(n1967), .CK(clk), .RN(n3368), .Q(
        \register_r[27][4] ), .QN(n294) );
  DFFRX1 \register_r_reg[27][3]  ( .D(n1966), .CK(clk), .RN(n3368), .Q(
        \register_r[27][3] ), .QN(n295) );
  DFFRX1 \register_r_reg[27][2]  ( .D(n1965), .CK(clk), .RN(n3368), .Q(
        \register_r[27][2] ), .QN(n296) );
  DFFRX1 \register_r_reg[27][1]  ( .D(n1964), .CK(clk), .RN(n3368), .Q(
        \register_r[27][1] ), .QN(n297) );
  DFFRX1 \register_r_reg[27][0]  ( .D(n1963), .CK(clk), .RN(n3368), .Q(
        \register_r[27][0] ), .QN(n298) );
  DFFRX1 \register_r_reg[23][23]  ( .D(n1858), .CK(clk), .RN(n3359), .Q(
        \register_r[23][23] ), .QN(n403) );
  DFFRX1 \register_r_reg[23][22]  ( .D(n1857), .CK(clk), .RN(n3359), .Q(
        \register_r[23][22] ), .QN(n404) );
  DFFRX1 \register_r_reg[23][21]  ( .D(n1856), .CK(clk), .RN(n3359), .Q(
        \register_r[23][21] ), .QN(n405) );
  DFFRX1 \register_r_reg[23][20]  ( .D(n1855), .CK(clk), .RN(n3359), .Q(
        \register_r[23][20] ), .QN(n406) );
  DFFRX1 \register_r_reg[23][19]  ( .D(n1854), .CK(clk), .RN(n3359), .Q(
        \register_r[23][19] ), .QN(n407) );
  DFFRX1 \register_r_reg[23][18]  ( .D(n1853), .CK(clk), .RN(n3359), .Q(
        \register_r[23][18] ), .QN(n408) );
  DFFRX1 \register_r_reg[23][17]  ( .D(n1852), .CK(clk), .RN(n3359), .Q(
        \register_r[23][17] ), .QN(n409) );
  DFFRX1 \register_r_reg[23][16]  ( .D(n1851), .CK(clk), .RN(n3359), .Q(
        \register_r[23][16] ), .QN(n410) );
  DFFRX1 \register_r_reg[23][15]  ( .D(n1850), .CK(clk), .RN(n3358), .Q(
        \register_r[23][15] ), .QN(n411) );
  DFFRX1 \register_r_reg[23][14]  ( .D(n1849), .CK(clk), .RN(n3358), .Q(
        \register_r[23][14] ), .QN(n412) );
  DFFRX1 \register_r_reg[23][13]  ( .D(n1848), .CK(clk), .RN(n3358), .Q(
        \register_r[23][13] ), .QN(n413) );
  DFFRX1 \register_r_reg[23][12]  ( .D(n1847), .CK(clk), .RN(n3358), .Q(
        \register_r[23][12] ), .QN(n414) );
  DFFRX1 \register_r_reg[23][11]  ( .D(n1846), .CK(clk), .RN(n3358), .Q(
        \register_r[23][11] ), .QN(n415) );
  DFFRX1 \register_r_reg[23][10]  ( .D(n1845), .CK(clk), .RN(n3358), .Q(
        \register_r[23][10] ), .QN(n416) );
  DFFRX1 \register_r_reg[23][9]  ( .D(n1844), .CK(clk), .RN(n3358), .Q(
        \register_r[23][9] ), .QN(n417) );
  DFFRX1 \register_r_reg[23][8]  ( .D(n1843), .CK(clk), .RN(n3358), .Q(
        \register_r[23][8] ), .QN(n418) );
  DFFRX1 \register_r_reg[23][7]  ( .D(n1842), .CK(clk), .RN(n3358), .Q(
        \register_r[23][7] ), .QN(n419) );
  DFFRX1 \register_r_reg[23][6]  ( .D(n1841), .CK(clk), .RN(n3358), .Q(
        \register_r[23][6] ), .QN(n420) );
  DFFRX1 \register_r_reg[23][5]  ( .D(n1840), .CK(clk), .RN(n3358), .Q(
        \register_r[23][5] ), .QN(n421) );
  DFFRX1 \register_r_reg[23][4]  ( .D(n1839), .CK(clk), .RN(n3358), .Q(
        \register_r[23][4] ), .QN(n422) );
  DFFRX1 \register_r_reg[23][3]  ( .D(n1838), .CK(clk), .RN(n3357), .Q(
        \register_r[23][3] ), .QN(n423) );
  DFFRX1 \register_r_reg[23][2]  ( .D(n1837), .CK(clk), .RN(n3357), .Q(
        \register_r[23][2] ), .QN(n424) );
  DFFRX1 \register_r_reg[23][1]  ( .D(n1836), .CK(clk), .RN(n3357), .Q(
        \register_r[23][1] ), .QN(n425) );
  DFFRX1 \register_r_reg[23][0]  ( .D(n1835), .CK(clk), .RN(n3357), .Q(
        \register_r[23][0] ), .QN(n426) );
  DFFRX1 \register_r_reg[19][23]  ( .D(n1730), .CK(clk), .RN(n3348), .Q(
        \register_r[19][23] ), .QN(n531) );
  DFFRX1 \register_r_reg[19][22]  ( .D(n1729), .CK(clk), .RN(n3348), .Q(
        \register_r[19][22] ), .QN(n532) );
  DFFRX1 \register_r_reg[19][21]  ( .D(n1728), .CK(clk), .RN(n3348), .Q(
        \register_r[19][21] ), .QN(n533) );
  DFFRX1 \register_r_reg[19][20]  ( .D(n1727), .CK(clk), .RN(n3348), .Q(
        \register_r[19][20] ), .QN(n534) );
  DFFRX1 \register_r_reg[19][19]  ( .D(n1726), .CK(clk), .RN(n3348), .Q(
        \register_r[19][19] ), .QN(n535) );
  DFFRX1 \register_r_reg[19][18]  ( .D(n1725), .CK(clk), .RN(n3348), .Q(
        \register_r[19][18] ), .QN(n536) );
  DFFRX1 \register_r_reg[19][17]  ( .D(n1724), .CK(clk), .RN(n3348), .Q(
        \register_r[19][17] ), .QN(n537) );
  DFFRX1 \register_r_reg[19][16]  ( .D(n1723), .CK(clk), .RN(n3348), .Q(
        \register_r[19][16] ), .QN(n538) );
  DFFRX1 \register_r_reg[19][15]  ( .D(n1722), .CK(clk), .RN(n3348), .Q(
        \register_r[19][15] ), .QN(n539) );
  DFFRX1 \register_r_reg[19][14]  ( .D(n1721), .CK(clk), .RN(n3348), .Q(
        \register_r[19][14] ), .QN(n540) );
  DFFRX1 \register_r_reg[19][13]  ( .D(n1720), .CK(clk), .RN(n3348), .Q(
        \register_r[19][13] ), .QN(n541) );
  DFFRX1 \register_r_reg[19][12]  ( .D(n1719), .CK(clk), .RN(n3348), .Q(
        \register_r[19][12] ), .QN(n542) );
  DFFRX1 \register_r_reg[19][11]  ( .D(n1718), .CK(clk), .RN(n3347), .Q(
        \register_r[19][11] ), .QN(n543) );
  DFFRX1 \register_r_reg[19][10]  ( .D(n1717), .CK(clk), .RN(n3347), .Q(
        \register_r[19][10] ), .QN(n544) );
  DFFRX1 \register_r_reg[19][9]  ( .D(n1716), .CK(clk), .RN(n3347), .Q(
        \register_r[19][9] ), .QN(n545) );
  DFFRX1 \register_r_reg[19][8]  ( .D(n1715), .CK(clk), .RN(n3347), .Q(
        \register_r[19][8] ), .QN(n546) );
  DFFRX1 \register_r_reg[19][7]  ( .D(n1714), .CK(clk), .RN(n3347), .Q(
        \register_r[19][7] ), .QN(n547) );
  DFFRX1 \register_r_reg[19][6]  ( .D(n1713), .CK(clk), .RN(n3347), .Q(
        \register_r[19][6] ), .QN(n548) );
  DFFRX1 \register_r_reg[19][5]  ( .D(n1712), .CK(clk), .RN(n3347), .Q(
        \register_r[19][5] ), .QN(n549) );
  DFFRX1 \register_r_reg[19][4]  ( .D(n1711), .CK(clk), .RN(n3347), .Q(
        \register_r[19][4] ), .QN(n550) );
  DFFRX1 \register_r_reg[19][3]  ( .D(n1710), .CK(clk), .RN(n3347), .Q(
        \register_r[19][3] ), .QN(n551) );
  DFFRX1 \register_r_reg[19][2]  ( .D(n1709), .CK(clk), .RN(n3347), .Q(
        \register_r[19][2] ), .QN(n552) );
  DFFRX1 \register_r_reg[19][1]  ( .D(n1708), .CK(clk), .RN(n3347), .Q(
        \register_r[19][1] ), .QN(n553) );
  DFFRX1 \register_r_reg[19][0]  ( .D(n1707), .CK(clk), .RN(n3347), .Q(
        \register_r[19][0] ), .QN(n554) );
  DFFRX1 \register_r_reg[15][31]  ( .D(n1610), .CK(clk), .RN(n3338), .Q(
        \register_r[15][31] ), .QN(n651) );
  DFFRX1 \register_r_reg[15][30]  ( .D(n1609), .CK(clk), .RN(n3338), .Q(
        \register_r[15][30] ), .QN(n652) );
  DFFRX1 \register_r_reg[15][29]  ( .D(n1608), .CK(clk), .RN(n3338), .Q(
        \register_r[15][29] ), .QN(n653) );
  DFFRX1 \register_r_reg[15][28]  ( .D(n1607), .CK(clk), .RN(n3338), .Q(
        \register_r[15][28] ), .QN(n654) );
  DFFRX1 \register_r_reg[15][27]  ( .D(n1606), .CK(clk), .RN(n3338), .Q(
        \register_r[15][27] ), .QN(n655) );
  DFFRX1 \register_r_reg[15][26]  ( .D(n1605), .CK(clk), .RN(n3338), .Q(
        \register_r[15][26] ), .QN(n656) );
  DFFRX1 \register_r_reg[15][25]  ( .D(n1604), .CK(clk), .RN(n3338), .Q(
        \register_r[15][25] ), .QN(n657) );
  DFFRX1 \register_r_reg[15][24]  ( .D(n1603), .CK(clk), .RN(n3338), .Q(
        \register_r[15][24] ), .QN(n658) );
  DFFRX1 \register_r_reg[15][23]  ( .D(n1602), .CK(clk), .RN(n3338), .Q(
        \register_r[15][23] ), .QN(n659) );
  DFFRX1 \register_r_reg[15][22]  ( .D(n1601), .CK(clk), .RN(n3338), .Q(
        \register_r[15][22] ), .QN(n660) );
  DFFRX1 \register_r_reg[15][21]  ( .D(n1600), .CK(clk), .RN(n3338), .Q(
        \register_r[15][21] ), .QN(n661) );
  DFFRX1 \register_r_reg[15][20]  ( .D(n1599), .CK(clk), .RN(n3338), .Q(
        \register_r[15][20] ), .QN(n662) );
  DFFRX1 \register_r_reg[15][19]  ( .D(n1598), .CK(clk), .RN(n3337), .Q(
        \register_r[15][19] ), .QN(n663) );
  DFFRX1 \register_r_reg[15][18]  ( .D(n1597), .CK(clk), .RN(n3337), .Q(
        \register_r[15][18] ), .QN(n664) );
  DFFRX1 \register_r_reg[15][17]  ( .D(n1596), .CK(clk), .RN(n3337), .Q(
        \register_r[15][17] ), .QN(n665) );
  DFFRX1 \register_r_reg[15][16]  ( .D(n1595), .CK(clk), .RN(n3337), .Q(
        \register_r[15][16] ), .QN(n666) );
  DFFRX1 \register_r_reg[15][15]  ( .D(n1594), .CK(clk), .RN(n3337), .Q(
        \register_r[15][15] ), .QN(n667) );
  DFFRX1 \register_r_reg[15][14]  ( .D(n1593), .CK(clk), .RN(n3337), .Q(
        \register_r[15][14] ), .QN(n668) );
  DFFRX1 \register_r_reg[15][13]  ( .D(n1592), .CK(clk), .RN(n3337), .Q(
        \register_r[15][13] ), .QN(n669) );
  DFFRX1 \register_r_reg[15][12]  ( .D(n1591), .CK(clk), .RN(n3337), .Q(
        \register_r[15][12] ), .QN(n670) );
  DFFRX1 \register_r_reg[15][11]  ( .D(n1590), .CK(clk), .RN(n3337), .Q(
        \register_r[15][11] ), .QN(n671) );
  DFFRX1 \register_r_reg[15][10]  ( .D(n1589), .CK(clk), .RN(n3337), .Q(
        \register_r[15][10] ), .QN(n672) );
  DFFRX1 \register_r_reg[15][9]  ( .D(n1588), .CK(clk), .RN(n3337), .Q(
        \register_r[15][9] ), .QN(n673) );
  DFFRX1 \register_r_reg[15][8]  ( .D(n1587), .CK(clk), .RN(n3337), .Q(
        \register_r[15][8] ), .QN(n674) );
  DFFRX1 \register_r_reg[15][7]  ( .D(n1586), .CK(clk), .RN(n3336), .Q(
        \register_r[15][7] ), .QN(n675) );
  DFFRX1 \register_r_reg[15][6]  ( .D(n1585), .CK(clk), .RN(n3336), .Q(
        \register_r[15][6] ), .QN(n676) );
  DFFRX1 \register_r_reg[15][5]  ( .D(n1584), .CK(clk), .RN(n3336), .Q(
        \register_r[15][5] ), .QN(n677) );
  DFFRX1 \register_r_reg[15][4]  ( .D(n1583), .CK(clk), .RN(n3336), .Q(
        \register_r[15][4] ), .QN(n678) );
  DFFRX1 \register_r_reg[15][3]  ( .D(n1582), .CK(clk), .RN(n3336), .Q(
        \register_r[15][3] ), .QN(n679) );
  DFFRX1 \register_r_reg[15][2]  ( .D(n1581), .CK(clk), .RN(n3336), .Q(
        \register_r[15][2] ), .QN(n680) );
  DFFRX1 \register_r_reg[15][1]  ( .D(n1580), .CK(clk), .RN(n3336), .Q(
        \register_r[15][1] ), .QN(n681) );
  DFFRX1 \register_r_reg[15][0]  ( .D(n1579), .CK(clk), .RN(n3336), .Q(
        \register_r[15][0] ), .QN(n682) );
  DFFRX1 \register_r_reg[11][31]  ( .D(n1482), .CK(clk), .RN(n3328), .Q(
        \register_r[11][31] ), .QN(n779) );
  DFFRX1 \register_r_reg[11][30]  ( .D(n1481), .CK(clk), .RN(n3328), .Q(
        \register_r[11][30] ), .QN(n780) );
  DFFRX1 \register_r_reg[11][29]  ( .D(n1480), .CK(clk), .RN(n3328), .Q(
        \register_r[11][29] ), .QN(n781) );
  DFFRX1 \register_r_reg[11][28]  ( .D(n1479), .CK(clk), .RN(n3328), .Q(
        \register_r[11][28] ), .QN(n782) );
  DFFRX1 \register_r_reg[11][27]  ( .D(n1478), .CK(clk), .RN(n3327), .Q(
        \register_r[11][27] ), .QN(n783) );
  DFFRX1 \register_r_reg[11][26]  ( .D(n1477), .CK(clk), .RN(n3327), .Q(
        \register_r[11][26] ), .QN(n784) );
  DFFRX1 \register_r_reg[11][25]  ( .D(n1476), .CK(clk), .RN(n3327), .Q(
        \register_r[11][25] ), .QN(n785) );
  DFFRX1 \register_r_reg[11][24]  ( .D(n1475), .CK(clk), .RN(n3327), .Q(
        \register_r[11][24] ), .QN(n786) );
  DFFRX1 \register_r_reg[11][23]  ( .D(n1474), .CK(clk), .RN(n3327), .Q(
        \register_r[11][23] ), .QN(n787) );
  DFFRX1 \register_r_reg[11][22]  ( .D(n1473), .CK(clk), .RN(n3327), .Q(
        \register_r[11][22] ), .QN(n788) );
  DFFRX1 \register_r_reg[11][21]  ( .D(n1472), .CK(clk), .RN(n3327), .Q(
        \register_r[11][21] ), .QN(n789) );
  DFFRX1 \register_r_reg[11][20]  ( .D(n1471), .CK(clk), .RN(n3327), .Q(
        \register_r[11][20] ), .QN(n790) );
  DFFRX1 \register_r_reg[11][19]  ( .D(n1470), .CK(clk), .RN(n3327), .Q(
        \register_r[11][19] ), .QN(n791) );
  DFFRX1 \register_r_reg[11][18]  ( .D(n1469), .CK(clk), .RN(n3327), .Q(
        \register_r[11][18] ), .QN(n792) );
  DFFRX1 \register_r_reg[11][17]  ( .D(n1468), .CK(clk), .RN(n3327), .Q(
        \register_r[11][17] ), .QN(n793) );
  DFFRX1 \register_r_reg[11][16]  ( .D(n1467), .CK(clk), .RN(n3327), .Q(
        \register_r[11][16] ), .QN(n794) );
  DFFRX1 \register_r_reg[11][15]  ( .D(n1466), .CK(clk), .RN(n3326), .Q(
        \register_r[11][15] ), .QN(n795) );
  DFFRX1 \register_r_reg[11][14]  ( .D(n1465), .CK(clk), .RN(n3326), .Q(
        \register_r[11][14] ), .QN(n796) );
  DFFRX1 \register_r_reg[11][13]  ( .D(n1464), .CK(clk), .RN(n3326), .Q(
        \register_r[11][13] ), .QN(n797) );
  DFFRX1 \register_r_reg[11][12]  ( .D(n1463), .CK(clk), .RN(n3326), .Q(
        \register_r[11][12] ), .QN(n798) );
  DFFRX1 \register_r_reg[11][11]  ( .D(n1462), .CK(clk), .RN(n3326), .Q(
        \register_r[11][11] ), .QN(n799) );
  DFFRX1 \register_r_reg[11][10]  ( .D(n1461), .CK(clk), .RN(n3326), .Q(
        \register_r[11][10] ), .QN(n800) );
  DFFRX1 \register_r_reg[11][9]  ( .D(n1460), .CK(clk), .RN(n3326), .Q(
        \register_r[11][9] ), .QN(n801) );
  DFFRX1 \register_r_reg[11][8]  ( .D(n1459), .CK(clk), .RN(n3326), .Q(
        \register_r[11][8] ), .QN(n802) );
  DFFRX1 \register_r_reg[11][7]  ( .D(n1458), .CK(clk), .RN(n3326), .Q(
        \register_r[11][7] ), .QN(n803) );
  DFFRX1 \register_r_reg[11][6]  ( .D(n1457), .CK(clk), .RN(n3326), .Q(
        \register_r[11][6] ), .QN(n804) );
  DFFRX1 \register_r_reg[11][5]  ( .D(n1456), .CK(clk), .RN(n3326), .Q(
        \register_r[11][5] ), .QN(n805) );
  DFFRX1 \register_r_reg[11][4]  ( .D(n1455), .CK(clk), .RN(n3326), .Q(
        \register_r[11][4] ), .QN(n806) );
  DFFRX1 \register_r_reg[11][3]  ( .D(n1454), .CK(clk), .RN(n3325), .Q(
        \register_r[11][3] ), .QN(n807) );
  DFFRX1 \register_r_reg[11][2]  ( .D(n1453), .CK(clk), .RN(n3325), .Q(
        \register_r[11][2] ), .QN(n808) );
  DFFRX1 \register_r_reg[11][1]  ( .D(n1452), .CK(clk), .RN(n3325), .Q(
        \register_r[11][1] ), .QN(n809) );
  DFFRX1 \register_r_reg[11][0]  ( .D(n1451), .CK(clk), .RN(n3325), .Q(
        \register_r[11][0] ), .QN(n810) );
  DFFRX1 \register_r_reg[7][31]  ( .D(n1354), .CK(clk), .RN(n3317), .Q(
        \register_r[7][31] ), .QN(n907) );
  DFFRX1 \register_r_reg[7][30]  ( .D(n1353), .CK(clk), .RN(n3317), .Q(
        \register_r[7][30] ), .QN(n908) );
  DFFRX1 \register_r_reg[7][29]  ( .D(n1352), .CK(clk), .RN(n3317), .Q(
        \register_r[7][29] ), .QN(n909) );
  DFFRX1 \register_r_reg[7][28]  ( .D(n1351), .CK(clk), .RN(n3317), .Q(
        \register_r[7][28] ), .QN(n910) );
  DFFRX1 \register_r_reg[7][27]  ( .D(n1350), .CK(clk), .RN(n3317), .Q(
        \register_r[7][27] ), .QN(n911) );
  DFFRX1 \register_r_reg[7][26]  ( .D(n1349), .CK(clk), .RN(n3317), .Q(
        \register_r[7][26] ), .QN(n912) );
  DFFRX1 \register_r_reg[7][25]  ( .D(n1348), .CK(clk), .RN(n3317), .Q(
        \register_r[7][25] ), .QN(n913) );
  DFFRX1 \register_r_reg[7][24]  ( .D(n1347), .CK(clk), .RN(n3317), .Q(
        \register_r[7][24] ), .QN(n914) );
  DFFRX1 \register_r_reg[7][23]  ( .D(n1346), .CK(clk), .RN(n3316), .Q(
        \register_r[7][23] ), .QN(n915) );
  DFFRX1 \register_r_reg[7][22]  ( .D(n1345), .CK(clk), .RN(n3316), .Q(
        \register_r[7][22] ), .QN(n916) );
  DFFRX1 \register_r_reg[7][21]  ( .D(n1344), .CK(clk), .RN(n3316), .Q(
        \register_r[7][21] ), .QN(n917) );
  DFFRX1 \register_r_reg[7][20]  ( .D(n1343), .CK(clk), .RN(n3316), .Q(
        \register_r[7][20] ), .QN(n918) );
  DFFRX1 \register_r_reg[7][19]  ( .D(n1342), .CK(clk), .RN(n3316), .Q(
        \register_r[7][19] ), .QN(n919) );
  DFFRX1 \register_r_reg[7][18]  ( .D(n1341), .CK(clk), .RN(n3316), .Q(
        \register_r[7][18] ), .QN(n920) );
  DFFRX1 \register_r_reg[7][17]  ( .D(n1340), .CK(clk), .RN(n3316), .Q(
        \register_r[7][17] ), .QN(n921) );
  DFFRX1 \register_r_reg[7][16]  ( .D(n1339), .CK(clk), .RN(n3316), .Q(
        \register_r[7][16] ), .QN(n922) );
  DFFRX1 \register_r_reg[7][15]  ( .D(n1338), .CK(clk), .RN(n3316), .Q(
        \register_r[7][15] ), .QN(n923) );
  DFFRX1 \register_r_reg[7][14]  ( .D(n1337), .CK(clk), .RN(n3316), .Q(
        \register_r[7][14] ), .QN(n924) );
  DFFRX1 \register_r_reg[7][13]  ( .D(n1336), .CK(clk), .RN(n3316), .Q(
        \register_r[7][13] ), .QN(n925) );
  DFFRX1 \register_r_reg[7][12]  ( .D(n1335), .CK(clk), .RN(n3316), .Q(
        \register_r[7][12] ), .QN(n926) );
  DFFRX1 \register_r_reg[7][11]  ( .D(n1334), .CK(clk), .RN(n3315), .Q(
        \register_r[7][11] ), .QN(n927) );
  DFFRX1 \register_r_reg[7][10]  ( .D(n1333), .CK(clk), .RN(n3315), .Q(
        \register_r[7][10] ), .QN(n928) );
  DFFRX1 \register_r_reg[7][9]  ( .D(n1332), .CK(clk), .RN(n3315), .Q(
        \register_r[7][9] ), .QN(n929) );
  DFFRX1 \register_r_reg[7][8]  ( .D(n1331), .CK(clk), .RN(n3315), .Q(
        \register_r[7][8] ), .QN(n930) );
  DFFRX1 \register_r_reg[7][7]  ( .D(n1330), .CK(clk), .RN(n3315), .Q(
        \register_r[7][7] ), .QN(n931) );
  DFFRX1 \register_r_reg[7][6]  ( .D(n1329), .CK(clk), .RN(n3315), .Q(
        \register_r[7][6] ), .QN(n932) );
  DFFRX1 \register_r_reg[7][5]  ( .D(n1328), .CK(clk), .RN(n3315), .Q(
        \register_r[7][5] ), .QN(n933) );
  DFFRX1 \register_r_reg[7][4]  ( .D(n1327), .CK(clk), .RN(n3315), .Q(
        \register_r[7][4] ), .QN(n934) );
  DFFRX1 \register_r_reg[7][3]  ( .D(n1326), .CK(clk), .RN(n3315), .Q(
        \register_r[7][3] ), .QN(n935) );
  DFFRX1 \register_r_reg[7][2]  ( .D(n1325), .CK(clk), .RN(n3315), .Q(
        \register_r[7][2] ), .QN(n936) );
  DFFRX1 \register_r_reg[7][1]  ( .D(n1324), .CK(clk), .RN(n3315), .Q(
        \register_r[7][1] ), .QN(n937) );
  DFFRX1 \register_r_reg[7][0]  ( .D(n1323), .CK(clk), .RN(n3315), .Q(
        \register_r[7][0] ), .QN(n938) );
  DFFRX1 \register_r_reg[29][31]  ( .D(n2058), .CK(clk), .RN(n3376), .Q(
        \register_r[29][31] ), .QN(n203) );
  DFFRX1 \register_r_reg[29][30]  ( .D(n2057), .CK(clk), .RN(n3376), .Q(
        \register_r[29][30] ), .QN(n204) );
  DFFRX1 \register_r_reg[29][29]  ( .D(n2056), .CK(clk), .RN(n3376), .Q(
        \register_r[29][29] ), .QN(n205) );
  DFFRX1 \register_r_reg[29][28]  ( .D(n2055), .CK(clk), .RN(n3376), .Q(
        \register_r[29][28] ), .QN(n206) );
  DFFRX1 \register_r_reg[29][27]  ( .D(n2054), .CK(clk), .RN(n3375), .Q(
        \register_r[29][27] ), .QN(n207) );
  DFFRX1 \register_r_reg[29][26]  ( .D(n2053), .CK(clk), .RN(n3375), .Q(
        \register_r[29][26] ), .QN(n208) );
  DFFRX1 \register_r_reg[29][25]  ( .D(n2052), .CK(clk), .RN(n3375), .Q(
        \register_r[29][25] ), .QN(n209) );
  DFFRX1 \register_r_reg[29][24]  ( .D(n2051), .CK(clk), .RN(n3375), .Q(
        \register_r[29][24] ), .QN(n210) );
  DFFRX1 \register_r_reg[29][23]  ( .D(n2050), .CK(clk), .RN(n3375), .Q(
        \register_r[29][23] ), .QN(n211) );
  DFFRX1 \register_r_reg[29][22]  ( .D(n2049), .CK(clk), .RN(n3375), .Q(
        \register_r[29][22] ), .QN(n212) );
  DFFRX1 \register_r_reg[29][21]  ( .D(n2048), .CK(clk), .RN(n3375), .Q(
        \register_r[29][21] ), .QN(n213) );
  DFFRX1 \register_r_reg[29][20]  ( .D(n2047), .CK(clk), .RN(n3375), .Q(
        \register_r[29][20] ), .QN(n214) );
  DFFRX1 \register_r_reg[29][19]  ( .D(n2046), .CK(clk), .RN(n3375), .Q(
        \register_r[29][19] ), .QN(n215) );
  DFFRX1 \register_r_reg[29][18]  ( .D(n2045), .CK(clk), .RN(n3375), .Q(
        \register_r[29][18] ), .QN(n216) );
  DFFRX1 \register_r_reg[29][17]  ( .D(n2044), .CK(clk), .RN(n3375), .Q(
        \register_r[29][17] ), .QN(n217) );
  DFFRX1 \register_r_reg[29][16]  ( .D(n2043), .CK(clk), .RN(n3375), .Q(
        \register_r[29][16] ), .QN(n218) );
  DFFRX1 \register_r_reg[29][15]  ( .D(n2042), .CK(clk), .RN(n3374), .Q(
        \register_r[29][15] ), .QN(n219) );
  DFFRX1 \register_r_reg[29][14]  ( .D(n2041), .CK(clk), .RN(n3374), .Q(
        \register_r[29][14] ), .QN(n220) );
  DFFRX1 \register_r_reg[29][13]  ( .D(n2040), .CK(clk), .RN(n3374), .Q(
        \register_r[29][13] ), .QN(n221) );
  DFFRX1 \register_r_reg[29][12]  ( .D(n2039), .CK(clk), .RN(n3374), .Q(
        \register_r[29][12] ), .QN(n222) );
  DFFRX1 \register_r_reg[29][11]  ( .D(n2038), .CK(clk), .RN(n3374), .Q(
        \register_r[29][11] ), .QN(n223) );
  DFFRX1 \register_r_reg[29][10]  ( .D(n2037), .CK(clk), .RN(n3374), .Q(
        \register_r[29][10] ), .QN(n224) );
  DFFRX1 \register_r_reg[29][9]  ( .D(n2036), .CK(clk), .RN(n3374), .Q(
        \register_r[29][9] ), .QN(n225) );
  DFFRX1 \register_r_reg[29][8]  ( .D(n2035), .CK(clk), .RN(n3374), .Q(
        \register_r[29][8] ), .QN(n226) );
  DFFRX1 \register_r_reg[29][7]  ( .D(n2034), .CK(clk), .RN(n3374), .Q(
        \register_r[29][7] ), .QN(n227) );
  DFFRX1 \register_r_reg[29][6]  ( .D(n2033), .CK(clk), .RN(n3374), .Q(
        \register_r[29][6] ), .QN(n228) );
  DFFRX1 \register_r_reg[29][5]  ( .D(n2032), .CK(clk), .RN(n3374), .Q(
        \register_r[29][5] ), .QN(n229) );
  DFFRX1 \register_r_reg[29][4]  ( .D(n2031), .CK(clk), .RN(n3374), .Q(
        \register_r[29][4] ), .QN(n230) );
  DFFRX1 \register_r_reg[29][3]  ( .D(n2030), .CK(clk), .RN(n3373), .Q(
        \register_r[29][3] ), .QN(n231) );
  DFFRX1 \register_r_reg[29][2]  ( .D(n2029), .CK(clk), .RN(n3373), .Q(
        \register_r[29][2] ), .QN(n232) );
  DFFRX1 \register_r_reg[29][1]  ( .D(n2028), .CK(clk), .RN(n3373), .Q(
        \register_r[29][1] ), .QN(n233) );
  DFFRX1 \register_r_reg[29][0]  ( .D(n2027), .CK(clk), .RN(n3373), .Q(
        \register_r[29][0] ), .QN(n234) );
  DFFRX1 \register_r_reg[25][31]  ( .D(n1930), .CK(clk), .RN(n3365), .Q(
        \register_r[25][31] ), .QN(n331) );
  DFFRX1 \register_r_reg[25][30]  ( .D(n1929), .CK(clk), .RN(n3365), .Q(
        \register_r[25][30] ), .QN(n332) );
  DFFRX1 \register_r_reg[25][29]  ( .D(n1928), .CK(clk), .RN(n3365), .Q(
        \register_r[25][29] ), .QN(n333) );
  DFFRX1 \register_r_reg[25][28]  ( .D(n1927), .CK(clk), .RN(n3365), .Q(
        \register_r[25][28] ), .QN(n334) );
  DFFRX1 \register_r_reg[25][27]  ( .D(n1926), .CK(clk), .RN(n3365), .Q(
        \register_r[25][27] ), .QN(n335) );
  DFFRX1 \register_r_reg[25][26]  ( .D(n1925), .CK(clk), .RN(n3365), .Q(
        \register_r[25][26] ), .QN(n336) );
  DFFRX1 \register_r_reg[25][25]  ( .D(n1924), .CK(clk), .RN(n3365), .Q(
        \register_r[25][25] ), .QN(n337) );
  DFFRX1 \register_r_reg[25][24]  ( .D(n1923), .CK(clk), .RN(n3365), .Q(
        \register_r[25][24] ), .QN(n338) );
  DFFRX1 \register_r_reg[25][23]  ( .D(n1922), .CK(clk), .RN(n3364), .Q(
        \register_r[25][23] ), .QN(n339) );
  DFFRX1 \register_r_reg[25][22]  ( .D(n1921), .CK(clk), .RN(n3364), .Q(
        \register_r[25][22] ), .QN(n340) );
  DFFRX1 \register_r_reg[25][21]  ( .D(n1920), .CK(clk), .RN(n3364), .Q(
        \register_r[25][21] ), .QN(n341) );
  DFFRX1 \register_r_reg[25][20]  ( .D(n1919), .CK(clk), .RN(n3364), .Q(
        \register_r[25][20] ), .QN(n342) );
  DFFRX1 \register_r_reg[25][19]  ( .D(n1918), .CK(clk), .RN(n3364), .Q(
        \register_r[25][19] ), .QN(n343) );
  DFFRX1 \register_r_reg[25][18]  ( .D(n1917), .CK(clk), .RN(n3364), .Q(
        \register_r[25][18] ), .QN(n344) );
  DFFRX1 \register_r_reg[25][17]  ( .D(n1916), .CK(clk), .RN(n3364), .Q(
        \register_r[25][17] ), .QN(n345) );
  DFFRX1 \register_r_reg[25][16]  ( .D(n1915), .CK(clk), .RN(n3364), .Q(
        \register_r[25][16] ), .QN(n346) );
  DFFRX1 \register_r_reg[25][15]  ( .D(n1914), .CK(clk), .RN(n3364), .Q(
        \register_r[25][15] ), .QN(n347) );
  DFFRX1 \register_r_reg[25][14]  ( .D(n1913), .CK(clk), .RN(n3364), .Q(
        \register_r[25][14] ), .QN(n348) );
  DFFRX1 \register_r_reg[25][13]  ( .D(n1912), .CK(clk), .RN(n3364), .Q(
        \register_r[25][13] ), .QN(n349) );
  DFFRX1 \register_r_reg[25][12]  ( .D(n1911), .CK(clk), .RN(n3364), .Q(
        \register_r[25][12] ), .QN(n350) );
  DFFRX1 \register_r_reg[25][11]  ( .D(n1910), .CK(clk), .RN(n3363), .Q(
        \register_r[25][11] ), .QN(n351) );
  DFFRX1 \register_r_reg[25][10]  ( .D(n1909), .CK(clk), .RN(n3363), .Q(
        \register_r[25][10] ), .QN(n352) );
  DFFRX1 \register_r_reg[25][9]  ( .D(n1908), .CK(clk), .RN(n3363), .Q(
        \register_r[25][9] ), .QN(n353) );
  DFFRX1 \register_r_reg[25][8]  ( .D(n1907), .CK(clk), .RN(n3363), .Q(
        \register_r[25][8] ), .QN(n354) );
  DFFRX1 \register_r_reg[25][7]  ( .D(n1906), .CK(clk), .RN(n3363), .Q(
        \register_r[25][7] ), .QN(n355) );
  DFFRX1 \register_r_reg[25][6]  ( .D(n1905), .CK(clk), .RN(n3363), .Q(
        \register_r[25][6] ), .QN(n356) );
  DFFRX1 \register_r_reg[25][5]  ( .D(n1904), .CK(clk), .RN(n3363), .Q(
        \register_r[25][5] ), .QN(n357) );
  DFFRX1 \register_r_reg[25][4]  ( .D(n1903), .CK(clk), .RN(n3363), .Q(
        \register_r[25][4] ), .QN(n358) );
  DFFRX1 \register_r_reg[25][3]  ( .D(n1902), .CK(clk), .RN(n3363), .Q(
        \register_r[25][3] ), .QN(n359) );
  DFFRX1 \register_r_reg[25][2]  ( .D(n1901), .CK(clk), .RN(n3363), .Q(
        \register_r[25][2] ), .QN(n360) );
  DFFRX1 \register_r_reg[25][1]  ( .D(n1900), .CK(clk), .RN(n3363), .Q(
        \register_r[25][1] ), .QN(n361) );
  DFFRX1 \register_r_reg[25][0]  ( .D(n1899), .CK(clk), .RN(n3363), .Q(
        \register_r[25][0] ), .QN(n362) );
  DFFRX1 \register_r_reg[21][23]  ( .D(n1794), .CK(clk), .RN(n3354), .Q(
        \register_r[21][23] ), .QN(n467) );
  DFFRX1 \register_r_reg[21][22]  ( .D(n1793), .CK(clk), .RN(n3354), .Q(
        \register_r[21][22] ), .QN(n468) );
  DFFRX1 \register_r_reg[21][21]  ( .D(n1792), .CK(clk), .RN(n3354), .Q(
        \register_r[21][21] ), .QN(n469) );
  DFFRX1 \register_r_reg[21][20]  ( .D(n1791), .CK(clk), .RN(n3354), .Q(
        \register_r[21][20] ), .QN(n470) );
  DFFRX1 \register_r_reg[21][19]  ( .D(n1790), .CK(clk), .RN(n3353), .Q(
        \register_r[21][19] ), .QN(n471) );
  DFFRX1 \register_r_reg[21][18]  ( .D(n1789), .CK(clk), .RN(n3353), .Q(
        \register_r[21][18] ), .QN(n472) );
  DFFRX1 \register_r_reg[21][17]  ( .D(n1788), .CK(clk), .RN(n3353), .Q(
        \register_r[21][17] ), .QN(n473) );
  DFFRX1 \register_r_reg[21][16]  ( .D(n1787), .CK(clk), .RN(n3353), .Q(
        \register_r[21][16] ), .QN(n474) );
  DFFRX1 \register_r_reg[21][15]  ( .D(n1786), .CK(clk), .RN(n3353), .Q(
        \register_r[21][15] ), .QN(n475) );
  DFFRX1 \register_r_reg[21][14]  ( .D(n1785), .CK(clk), .RN(n3353), .Q(
        \register_r[21][14] ), .QN(n476) );
  DFFRX1 \register_r_reg[21][13]  ( .D(n1784), .CK(clk), .RN(n3353), .Q(
        \register_r[21][13] ), .QN(n477) );
  DFFRX1 \register_r_reg[21][12]  ( .D(n1783), .CK(clk), .RN(n3353), .Q(
        \register_r[21][12] ), .QN(n478) );
  DFFRX1 \register_r_reg[21][11]  ( .D(n1782), .CK(clk), .RN(n3353), .Q(
        \register_r[21][11] ), .QN(n479) );
  DFFRX1 \register_r_reg[21][10]  ( .D(n1781), .CK(clk), .RN(n3353), .Q(
        \register_r[21][10] ), .QN(n480) );
  DFFRX1 \register_r_reg[21][9]  ( .D(n1780), .CK(clk), .RN(n3353), .Q(
        \register_r[21][9] ), .QN(n481) );
  DFFRX1 \register_r_reg[21][8]  ( .D(n1779), .CK(clk), .RN(n3353), .Q(
        \register_r[21][8] ), .QN(n482) );
  DFFRX1 \register_r_reg[21][7]  ( .D(n1778), .CK(clk), .RN(n3352), .Q(
        \register_r[21][7] ), .QN(n483) );
  DFFRX1 \register_r_reg[21][6]  ( .D(n1777), .CK(clk), .RN(n3352), .Q(
        \register_r[21][6] ), .QN(n484) );
  DFFRX1 \register_r_reg[21][5]  ( .D(n1776), .CK(clk), .RN(n3352), .Q(
        \register_r[21][5] ), .QN(n485) );
  DFFRX1 \register_r_reg[21][4]  ( .D(n1775), .CK(clk), .RN(n3352), .Q(
        \register_r[21][4] ), .QN(n486) );
  DFFRX1 \register_r_reg[21][3]  ( .D(n1774), .CK(clk), .RN(n3352), .Q(
        \register_r[21][3] ), .QN(n487) );
  DFFRX1 \register_r_reg[21][2]  ( .D(n1773), .CK(clk), .RN(n3352), .Q(
        \register_r[21][2] ), .QN(n488) );
  DFFRX1 \register_r_reg[21][1]  ( .D(n1772), .CK(clk), .RN(n3352), .Q(
        \register_r[21][1] ), .QN(n489) );
  DFFRX1 \register_r_reg[21][0]  ( .D(n1771), .CK(clk), .RN(n3352), .Q(
        \register_r[21][0] ), .QN(n490) );
  DFFRX1 \register_r_reg[17][28]  ( .D(n1671), .CK(clk), .RN(n3344), .Q(
        \register_r[17][28] ), .QN(n590) );
  DFFRX1 \register_r_reg[17][27]  ( .D(n1670), .CK(clk), .RN(n3343), .Q(
        \register_r[17][27] ), .QN(n591) );
  DFFRX1 \register_r_reg[17][26]  ( .D(n1669), .CK(clk), .RN(n3343), .Q(
        \register_r[17][26] ), .QN(n592) );
  DFFRX1 \register_r_reg[17][25]  ( .D(n1668), .CK(clk), .RN(n3343), .Q(
        \register_r[17][25] ), .QN(n593) );
  DFFRX1 \register_r_reg[17][24]  ( .D(n1667), .CK(clk), .RN(n3343), .Q(
        \register_r[17][24] ), .QN(n594) );
  DFFRX1 \register_r_reg[17][23]  ( .D(n1666), .CK(clk), .RN(n3343), .Q(
        \register_r[17][23] ), .QN(n595) );
  DFFRX1 \register_r_reg[17][22]  ( .D(n1665), .CK(clk), .RN(n3343), .Q(
        \register_r[17][22] ), .QN(n596) );
  DFFRX1 \register_r_reg[17][21]  ( .D(n1664), .CK(clk), .RN(n3343), .Q(
        \register_r[17][21] ), .QN(n597) );
  DFFRX1 \register_r_reg[17][20]  ( .D(n1663), .CK(clk), .RN(n3343), .Q(
        \register_r[17][20] ), .QN(n598) );
  DFFRX1 \register_r_reg[17][19]  ( .D(n1662), .CK(clk), .RN(n3343), .Q(
        \register_r[17][19] ), .QN(n599) );
  DFFRX1 \register_r_reg[17][18]  ( .D(n1661), .CK(clk), .RN(n3343), .Q(
        \register_r[17][18] ), .QN(n600) );
  DFFRX1 \register_r_reg[17][17]  ( .D(n1660), .CK(clk), .RN(n3343), .Q(
        \register_r[17][17] ), .QN(n601) );
  DFFRX1 \register_r_reg[17][16]  ( .D(n1659), .CK(clk), .RN(n3343), .Q(
        \register_r[17][16] ), .QN(n602) );
  DFFRX1 \register_r_reg[17][15]  ( .D(n1658), .CK(clk), .RN(n3342), .Q(
        \register_r[17][15] ), .QN(n603) );
  DFFRX1 \register_r_reg[17][14]  ( .D(n1657), .CK(clk), .RN(n3342), .Q(
        \register_r[17][14] ), .QN(n604) );
  DFFRX1 \register_r_reg[17][13]  ( .D(n1656), .CK(clk), .RN(n3342), .Q(
        \register_r[17][13] ), .QN(n605) );
  DFFRX1 \register_r_reg[17][12]  ( .D(n1655), .CK(clk), .RN(n3342), .Q(
        \register_r[17][12] ), .QN(n606) );
  DFFRX1 \register_r_reg[17][11]  ( .D(n1654), .CK(clk), .RN(n3342), .Q(
        \register_r[17][11] ), .QN(n607) );
  DFFRX1 \register_r_reg[17][10]  ( .D(n1653), .CK(clk), .RN(n3342), .Q(
        \register_r[17][10] ), .QN(n608) );
  DFFRX1 \register_r_reg[17][9]  ( .D(n1652), .CK(clk), .RN(n3342), .Q(
        \register_r[17][9] ), .QN(n609) );
  DFFRX1 \register_r_reg[17][8]  ( .D(n1651), .CK(clk), .RN(n3342), .Q(
        \register_r[17][8] ), .QN(n610) );
  DFFRX1 \register_r_reg[17][7]  ( .D(n1650), .CK(clk), .RN(n3342), .Q(
        \register_r[17][7] ), .QN(n611) );
  DFFRX1 \register_r_reg[17][6]  ( .D(n1649), .CK(clk), .RN(n3342), .Q(
        \register_r[17][6] ), .QN(n612) );
  DFFRX1 \register_r_reg[17][5]  ( .D(n1648), .CK(clk), .RN(n3342), .Q(
        \register_r[17][5] ), .QN(n613) );
  DFFRX1 \register_r_reg[17][4]  ( .D(n1647), .CK(clk), .RN(n3342), .Q(
        \register_r[17][4] ), .QN(n614) );
  DFFRX1 \register_r_reg[17][3]  ( .D(n1646), .CK(clk), .RN(n3341), .Q(
        \register_r[17][3] ), .QN(n615) );
  DFFRX1 \register_r_reg[17][2]  ( .D(n1645), .CK(clk), .RN(n3341), .Q(
        \register_r[17][2] ), .QN(n616) );
  DFFRX1 \register_r_reg[17][1]  ( .D(n1644), .CK(clk), .RN(n3341), .Q(
        \register_r[17][1] ), .QN(n617) );
  DFFRX1 \register_r_reg[17][0]  ( .D(n1643), .CK(clk), .RN(n3341), .Q(
        \register_r[17][0] ), .QN(n618) );
  DFFRX1 \register_r_reg[13][31]  ( .D(n1546), .CK(clk), .RN(n3333), .Q(
        r_13[31]), .QN(n715) );
  DFFRX1 \register_r_reg[13][30]  ( .D(n1545), .CK(clk), .RN(n3333), .Q(
        r_13[30]), .QN(n716) );
  DFFRX1 \register_r_reg[13][29]  ( .D(n1544), .CK(clk), .RN(n3333), .Q(
        r_13[29]), .QN(n717) );
  DFFRX1 \register_r_reg[13][28]  ( .D(n1543), .CK(clk), .RN(n3333), .Q(
        r_13[28]), .QN(n718) );
  DFFRX1 \register_r_reg[13][27]  ( .D(n1542), .CK(clk), .RN(n3333), .Q(
        r_13[27]), .QN(n719) );
  DFFRX1 \register_r_reg[13][26]  ( .D(n1541), .CK(clk), .RN(n3333), .Q(
        r_13[26]), .QN(n720) );
  DFFRX1 \register_r_reg[13][25]  ( .D(n1540), .CK(clk), .RN(n3333), .Q(
        r_13[25]), .QN(n721) );
  DFFRX1 \register_r_reg[13][24]  ( .D(n1539), .CK(clk), .RN(n3333), .Q(
        r_13[24]), .QN(n722) );
  DFFRX1 \register_r_reg[13][23]  ( .D(n1538), .CK(clk), .RN(n3332), .Q(
        r_13[23]), .QN(n723) );
  DFFRX1 \register_r_reg[13][22]  ( .D(n1537), .CK(clk), .RN(n3332), .Q(
        r_13[22]), .QN(n724) );
  DFFRX1 \register_r_reg[13][21]  ( .D(n1536), .CK(clk), .RN(n3332), .Q(
        r_13[21]), .QN(n725) );
  DFFRX1 \register_r_reg[13][20]  ( .D(n1535), .CK(clk), .RN(n3332), .Q(
        r_13[20]), .QN(n726) );
  DFFRX1 \register_r_reg[13][19]  ( .D(n1534), .CK(clk), .RN(n3332), .Q(
        r_13[19]), .QN(n727) );
  DFFRX1 \register_r_reg[13][18]  ( .D(n1533), .CK(clk), .RN(n3332), .Q(
        r_13[18]), .QN(n728) );
  DFFRX1 \register_r_reg[13][17]  ( .D(n1532), .CK(clk), .RN(n3332), .Q(
        r_13[17]), .QN(n729) );
  DFFRX1 \register_r_reg[13][16]  ( .D(n1531), .CK(clk), .RN(n3332), .Q(
        r_13[16]), .QN(n730) );
  DFFRX1 \register_r_reg[13][15]  ( .D(n1530), .CK(clk), .RN(n3332), .Q(
        r_13[15]), .QN(n731) );
  DFFRX1 \register_r_reg[13][14]  ( .D(n1529), .CK(clk), .RN(n3332), .Q(
        r_13[14]), .QN(n732) );
  DFFRX1 \register_r_reg[13][13]  ( .D(n1528), .CK(clk), .RN(n3332), .Q(
        r_13[13]), .QN(n733) );
  DFFRX1 \register_r_reg[13][12]  ( .D(n1527), .CK(clk), .RN(n3332), .Q(
        r_13[12]), .QN(n734) );
  DFFRX1 \register_r_reg[13][11]  ( .D(n1526), .CK(clk), .RN(n3331), .Q(
        r_13[11]), .QN(n735) );
  DFFRX1 \register_r_reg[13][10]  ( .D(n1525), .CK(clk), .RN(n3331), .Q(
        r_13[10]), .QN(n736) );
  DFFRX1 \register_r_reg[13][9]  ( .D(n1524), .CK(clk), .RN(n3331), .Q(r_13[9]), .QN(n737) );
  DFFRX1 \register_r_reg[13][8]  ( .D(n1523), .CK(clk), .RN(n3331), .Q(r_13[8]), .QN(n738) );
  DFFRX1 \register_r_reg[13][7]  ( .D(n1522), .CK(clk), .RN(n3331), .Q(r_13[7]), .QN(n739) );
  DFFRX1 \register_r_reg[13][6]  ( .D(n1521), .CK(clk), .RN(n3331), .Q(r_13[6]), .QN(n740) );
  DFFRX1 \register_r_reg[13][5]  ( .D(n1520), .CK(clk), .RN(n3331), .Q(r_13[5]), .QN(n741) );
  DFFRX1 \register_r_reg[13][4]  ( .D(n1519), .CK(clk), .RN(n3331), .Q(r_13[4]), .QN(n742) );
  DFFRX1 \register_r_reg[13][3]  ( .D(n1518), .CK(clk), .RN(n3331), .Q(r_13[3]), .QN(n743) );
  DFFRX1 \register_r_reg[13][2]  ( .D(n1517), .CK(clk), .RN(n3331), .Q(r_13[2]), .QN(n744) );
  DFFRX1 \register_r_reg[13][1]  ( .D(n1516), .CK(clk), .RN(n3331), .Q(r_13[1]), .QN(n745) );
  DFFRX1 \register_r_reg[13][0]  ( .D(n1515), .CK(clk), .RN(n3331), .Q(r_13[0]), .QN(n746) );
  DFFRX1 \register_r_reg[9][31]  ( .D(n1418), .CK(clk), .RN(n3322), .Q(
        \register_r[9][31] ), .QN(n843) );
  DFFRX1 \register_r_reg[9][30]  ( .D(n1417), .CK(clk), .RN(n3322), .Q(
        \register_r[9][30] ), .QN(n844) );
  DFFRX1 \register_r_reg[9][29]  ( .D(n1416), .CK(clk), .RN(n3322), .Q(
        \register_r[9][29] ), .QN(n845) );
  DFFRX1 \register_r_reg[9][28]  ( .D(n1415), .CK(clk), .RN(n3322), .Q(
        \register_r[9][28] ), .QN(n846) );
  DFFRX1 \register_r_reg[9][27]  ( .D(n1414), .CK(clk), .RN(n3322), .Q(
        \register_r[9][27] ), .QN(n847) );
  DFFRX1 \register_r_reg[9][26]  ( .D(n1413), .CK(clk), .RN(n3322), .Q(
        \register_r[9][26] ), .QN(n848) );
  DFFRX1 \register_r_reg[9][25]  ( .D(n1412), .CK(clk), .RN(n3322), .Q(
        \register_r[9][25] ), .QN(n849) );
  DFFRX1 \register_r_reg[9][24]  ( .D(n1411), .CK(clk), .RN(n3322), .Q(
        \register_r[9][24] ), .QN(n850) );
  DFFRX1 \register_r_reg[9][23]  ( .D(n1410), .CK(clk), .RN(n3322), .Q(
        \register_r[9][23] ), .QN(n851) );
  DFFRX1 \register_r_reg[9][22]  ( .D(n1409), .CK(clk), .RN(n3322), .Q(
        \register_r[9][22] ), .QN(n852) );
  DFFRX1 \register_r_reg[9][21]  ( .D(n1408), .CK(clk), .RN(n3322), .Q(
        \register_r[9][21] ), .QN(n853) );
  DFFRX1 \register_r_reg[9][20]  ( .D(n1407), .CK(clk), .RN(n3322), .Q(
        \register_r[9][20] ), .QN(n854) );
  DFFRX1 \register_r_reg[9][19]  ( .D(n1406), .CK(clk), .RN(n3321), .Q(
        \register_r[9][19] ), .QN(n855) );
  DFFRX1 \register_r_reg[9][18]  ( .D(n1405), .CK(clk), .RN(n3321), .Q(
        \register_r[9][18] ), .QN(n856) );
  DFFRX1 \register_r_reg[9][17]  ( .D(n1404), .CK(clk), .RN(n3321), .Q(
        \register_r[9][17] ), .QN(n857) );
  DFFRX1 \register_r_reg[9][16]  ( .D(n1403), .CK(clk), .RN(n3321), .Q(
        \register_r[9][16] ), .QN(n858) );
  DFFRX1 \register_r_reg[9][15]  ( .D(n1402), .CK(clk), .RN(n3321), .Q(
        \register_r[9][15] ), .QN(n859) );
  DFFRX1 \register_r_reg[9][14]  ( .D(n1401), .CK(clk), .RN(n3321), .Q(
        \register_r[9][14] ), .QN(n860) );
  DFFRX1 \register_r_reg[9][13]  ( .D(n1400), .CK(clk), .RN(n3321), .Q(
        \register_r[9][13] ), .QN(n861) );
  DFFRX1 \register_r_reg[9][12]  ( .D(n1399), .CK(clk), .RN(n3321), .Q(
        \register_r[9][12] ), .QN(n862) );
  DFFRX1 \register_r_reg[9][11]  ( .D(n1398), .CK(clk), .RN(n3321), .Q(
        \register_r[9][11] ), .QN(n863) );
  DFFRX1 \register_r_reg[9][10]  ( .D(n1397), .CK(clk), .RN(n3321), .Q(
        \register_r[9][10] ), .QN(n864) );
  DFFRX1 \register_r_reg[9][9]  ( .D(n1396), .CK(clk), .RN(n3321), .Q(
        \register_r[9][9] ), .QN(n865) );
  DFFRX1 \register_r_reg[9][8]  ( .D(n1395), .CK(clk), .RN(n3321), .Q(
        \register_r[9][8] ), .QN(n866) );
  DFFRX1 \register_r_reg[9][7]  ( .D(n1394), .CK(clk), .RN(n3320), .Q(
        \register_r[9][7] ), .QN(n867) );
  DFFRX1 \register_r_reg[9][6]  ( .D(n1393), .CK(clk), .RN(n3320), .Q(
        \register_r[9][6] ), .QN(n868) );
  DFFRX1 \register_r_reg[9][5]  ( .D(n1392), .CK(clk), .RN(n3320), .Q(
        \register_r[9][5] ), .QN(n869) );
  DFFRX1 \register_r_reg[9][4]  ( .D(n1391), .CK(clk), .RN(n3320), .Q(
        \register_r[9][4] ), .QN(n870) );
  DFFRX1 \register_r_reg[9][3]  ( .D(n1390), .CK(clk), .RN(n3320), .Q(
        \register_r[9][3] ), .QN(n871) );
  DFFRX1 \register_r_reg[9][2]  ( .D(n1389), .CK(clk), .RN(n3320), .Q(
        \register_r[9][2] ), .QN(n872) );
  DFFRX1 \register_r_reg[9][1]  ( .D(n1388), .CK(clk), .RN(n3320), .Q(
        \register_r[9][1] ), .QN(n873) );
  DFFRX1 \register_r_reg[9][0]  ( .D(n1387), .CK(clk), .RN(n3320), .Q(
        \register_r[9][0] ), .QN(n874) );
  DFFRX1 \register_r_reg[5][31]  ( .D(n1290), .CK(clk), .RN(n3312), .Q(
        \register_r[5][31] ), .QN(n971) );
  DFFRX1 \register_r_reg[5][30]  ( .D(n1289), .CK(clk), .RN(n3312), .Q(
        \register_r[5][30] ), .QN(n972) );
  DFFRX1 \register_r_reg[5][29]  ( .D(n1288), .CK(clk), .RN(n3312), .Q(
        \register_r[5][29] ), .QN(n973) );
  DFFRX1 \register_r_reg[5][28]  ( .D(n1287), .CK(clk), .RN(n3312), .Q(
        \register_r[5][28] ), .QN(n974) );
  DFFRX1 \register_r_reg[5][27]  ( .D(n1286), .CK(clk), .RN(n3311), .Q(
        \register_r[5][27] ), .QN(n975) );
  DFFRX1 \register_r_reg[5][26]  ( .D(n1285), .CK(clk), .RN(n3311), .Q(
        \register_r[5][26] ), .QN(n976) );
  DFFRX1 \register_r_reg[5][25]  ( .D(n1284), .CK(clk), .RN(n3311), .Q(
        \register_r[5][25] ), .QN(n977) );
  DFFRX1 \register_r_reg[5][24]  ( .D(n1283), .CK(clk), .RN(n3311), .Q(
        \register_r[5][24] ), .QN(n978) );
  DFFRX1 \register_r_reg[5][23]  ( .D(n1282), .CK(clk), .RN(n3311), .Q(
        \register_r[5][23] ), .QN(n979) );
  DFFRX1 \register_r_reg[5][22]  ( .D(n1281), .CK(clk), .RN(n3311), .Q(
        \register_r[5][22] ), .QN(n980) );
  DFFRX1 \register_r_reg[5][21]  ( .D(n1280), .CK(clk), .RN(n3311), .Q(
        \register_r[5][21] ), .QN(n981) );
  DFFRX1 \register_r_reg[5][20]  ( .D(n1279), .CK(clk), .RN(n3311), .Q(
        \register_r[5][20] ), .QN(n982) );
  DFFRX1 \register_r_reg[5][19]  ( .D(n1278), .CK(clk), .RN(n3311), .Q(
        \register_r[5][19] ), .QN(n983) );
  DFFRX1 \register_r_reg[5][18]  ( .D(n1277), .CK(clk), .RN(n3311), .Q(
        \register_r[5][18] ), .QN(n984) );
  DFFRX1 \register_r_reg[5][17]  ( .D(n1276), .CK(clk), .RN(n3311), .Q(
        \register_r[5][17] ), .QN(n985) );
  DFFRX1 \register_r_reg[5][16]  ( .D(n1275), .CK(clk), .RN(n3311), .Q(
        \register_r[5][16] ), .QN(n986) );
  DFFRX1 \register_r_reg[5][15]  ( .D(n1274), .CK(clk), .RN(n3310), .Q(
        \register_r[5][15] ), .QN(n987) );
  DFFRX1 \register_r_reg[5][14]  ( .D(n1273), .CK(clk), .RN(n3310), .Q(
        \register_r[5][14] ), .QN(n988) );
  DFFRX1 \register_r_reg[5][13]  ( .D(n1272), .CK(clk), .RN(n3310), .Q(
        \register_r[5][13] ), .QN(n989) );
  DFFRX1 \register_r_reg[5][12]  ( .D(n1271), .CK(clk), .RN(n3310), .Q(
        \register_r[5][12] ), .QN(n990) );
  DFFRX1 \register_r_reg[5][11]  ( .D(n1270), .CK(clk), .RN(n3310), .Q(
        \register_r[5][11] ), .QN(n991) );
  DFFRX1 \register_r_reg[5][10]  ( .D(n1269), .CK(clk), .RN(n3310), .Q(
        \register_r[5][10] ), .QN(n992) );
  DFFRX1 \register_r_reg[5][9]  ( .D(n1268), .CK(clk), .RN(n3310), .Q(
        \register_r[5][9] ), .QN(n993) );
  DFFRX1 \register_r_reg[5][8]  ( .D(n1267), .CK(clk), .RN(n3310), .Q(
        \register_r[5][8] ), .QN(n994) );
  DFFRX1 \register_r_reg[5][7]  ( .D(n1266), .CK(clk), .RN(n3310), .Q(
        \register_r[5][7] ), .QN(n995) );
  DFFRX1 \register_r_reg[5][6]  ( .D(n1265), .CK(clk), .RN(n3310), .Q(
        \register_r[5][6] ), .QN(n996) );
  DFFRX1 \register_r_reg[5][5]  ( .D(n1264), .CK(clk), .RN(n3310), .Q(
        \register_r[5][5] ), .QN(n997) );
  DFFRX1 \register_r_reg[5][4]  ( .D(n1263), .CK(clk), .RN(n3310), .Q(
        \register_r[5][4] ), .QN(n998) );
  DFFRX1 \register_r_reg[5][3]  ( .D(n1262), .CK(clk), .RN(n3309), .Q(
        \register_r[5][3] ), .QN(n999) );
  DFFRX1 \register_r_reg[5][2]  ( .D(n1261), .CK(clk), .RN(n3309), .Q(
        \register_r[5][2] ), .QN(n1000) );
  DFFRX1 \register_r_reg[5][1]  ( .D(n1260), .CK(clk), .RN(n3309), .Q(
        \register_r[5][1] ), .QN(n1001) );
  DFFRX1 \register_r_reg[5][0]  ( .D(n1259), .CK(clk), .RN(n3309), .Q(
        \register_r[5][0] ), .QN(n1002) );
  DFFRX1 \register_r_reg[28][31]  ( .D(n2026), .CK(clk), .RN(n3373), .Q(
        \register_r[28][31] ), .QN(n235) );
  DFFRX1 \register_r_reg[28][30]  ( .D(n2025), .CK(clk), .RN(n3373), .Q(
        \register_r[28][30] ), .QN(n236) );
  DFFRX1 \register_r_reg[28][29]  ( .D(n2024), .CK(clk), .RN(n3373), .Q(
        \register_r[28][29] ), .QN(n237) );
  DFFRX1 \register_r_reg[28][28]  ( .D(n2023), .CK(clk), .RN(n3373), .Q(
        \register_r[28][28] ), .QN(n238) );
  DFFRX1 \register_r_reg[28][27]  ( .D(n2022), .CK(clk), .RN(n3373), .Q(
        \register_r[28][27] ), .QN(n239) );
  DFFRX1 \register_r_reg[28][26]  ( .D(n2021), .CK(clk), .RN(n3373), .Q(
        \register_r[28][26] ), .QN(n240) );
  DFFRX1 \register_r_reg[28][25]  ( .D(n2020), .CK(clk), .RN(n3373), .Q(
        \register_r[28][25] ), .QN(n241) );
  DFFRX1 \register_r_reg[28][24]  ( .D(n2019), .CK(clk), .RN(n3373), .Q(
        \register_r[28][24] ), .QN(n242) );
  DFFRX1 \register_r_reg[28][23]  ( .D(n2018), .CK(clk), .RN(n3372), .Q(
        \register_r[28][23] ), .QN(n243) );
  DFFRX1 \register_r_reg[28][22]  ( .D(n2017), .CK(clk), .RN(n3372), .Q(
        \register_r[28][22] ), .QN(n244) );
  DFFRX1 \register_r_reg[28][21]  ( .D(n2016), .CK(clk), .RN(n3372), .Q(
        \register_r[28][21] ), .QN(n245) );
  DFFRX1 \register_r_reg[28][20]  ( .D(n2015), .CK(clk), .RN(n3372), .Q(
        \register_r[28][20] ), .QN(n246) );
  DFFRX1 \register_r_reg[28][19]  ( .D(n2014), .CK(clk), .RN(n3372), .Q(
        \register_r[28][19] ), .QN(n247) );
  DFFRX1 \register_r_reg[28][18]  ( .D(n2013), .CK(clk), .RN(n3372), .Q(
        \register_r[28][18] ), .QN(n248) );
  DFFRX1 \register_r_reg[28][17]  ( .D(n2012), .CK(clk), .RN(n3372), .Q(
        \register_r[28][17] ), .QN(n249) );
  DFFRX1 \register_r_reg[28][16]  ( .D(n2011), .CK(clk), .RN(n3372), .Q(
        \register_r[28][16] ), .QN(n250) );
  DFFRX1 \register_r_reg[28][15]  ( .D(n2010), .CK(clk), .RN(n3372), .Q(
        \register_r[28][15] ), .QN(n251) );
  DFFRX1 \register_r_reg[28][14]  ( .D(n2009), .CK(clk), .RN(n3372), .Q(
        \register_r[28][14] ), .QN(n252) );
  DFFRX1 \register_r_reg[28][13]  ( .D(n2008), .CK(clk), .RN(n3372), .Q(
        \register_r[28][13] ), .QN(n253) );
  DFFRX1 \register_r_reg[28][12]  ( .D(n2007), .CK(clk), .RN(n3372), .Q(
        \register_r[28][12] ), .QN(n254) );
  DFFRX1 \register_r_reg[28][11]  ( .D(n2006), .CK(clk), .RN(n3371), .Q(
        \register_r[28][11] ), .QN(n255) );
  DFFRX1 \register_r_reg[28][10]  ( .D(n2005), .CK(clk), .RN(n3371), .Q(
        \register_r[28][10] ), .QN(n256) );
  DFFRX1 \register_r_reg[28][9]  ( .D(n2004), .CK(clk), .RN(n3371), .Q(
        \register_r[28][9] ), .QN(n257) );
  DFFRX1 \register_r_reg[28][8]  ( .D(n2003), .CK(clk), .RN(n3371), .Q(
        \register_r[28][8] ), .QN(n258) );
  DFFRX1 \register_r_reg[28][7]  ( .D(n2002), .CK(clk), .RN(n3371), .Q(
        \register_r[28][7] ), .QN(n259) );
  DFFRX1 \register_r_reg[28][6]  ( .D(n2001), .CK(clk), .RN(n3371), .Q(
        \register_r[28][6] ), .QN(n260) );
  DFFRX1 \register_r_reg[28][5]  ( .D(n2000), .CK(clk), .RN(n3371), .Q(
        \register_r[28][5] ), .QN(n261) );
  DFFRX1 \register_r_reg[28][4]  ( .D(n1999), .CK(clk), .RN(n3371), .Q(
        \register_r[28][4] ), .QN(n262) );
  DFFRX1 \register_r_reg[28][3]  ( .D(n1998), .CK(clk), .RN(n3371), .Q(
        \register_r[28][3] ), .QN(n263) );
  DFFRX1 \register_r_reg[28][2]  ( .D(n1997), .CK(clk), .RN(n3371), .Q(
        \register_r[28][2] ), .QN(n264) );
  DFFRX1 \register_r_reg[28][1]  ( .D(n1996), .CK(clk), .RN(n3371), .Q(
        \register_r[28][1] ), .QN(n265) );
  DFFRX1 \register_r_reg[28][0]  ( .D(n1995), .CK(clk), .RN(n3371), .Q(
        \register_r[28][0] ), .QN(n266) );
  DFFRX1 \register_r_reg[24][31]  ( .D(n1898), .CK(clk), .RN(n3362), .Q(
        \register_r[24][31] ), .QN(n363) );
  DFFRX1 \register_r_reg[24][30]  ( .D(n1897), .CK(clk), .RN(n3362), .Q(
        \register_r[24][30] ), .QN(n364) );
  DFFRX1 \register_r_reg[24][29]  ( .D(n1896), .CK(clk), .RN(n3362), .Q(
        \register_r[24][29] ), .QN(n365) );
  DFFRX1 \register_r_reg[24][28]  ( .D(n1895), .CK(clk), .RN(n3362), .Q(
        \register_r[24][28] ), .QN(n366) );
  DFFRX1 \register_r_reg[24][27]  ( .D(n1894), .CK(clk), .RN(n3362), .Q(
        \register_r[24][27] ), .QN(n367) );
  DFFRX1 \register_r_reg[24][26]  ( .D(n1893), .CK(clk), .RN(n3362), .Q(
        \register_r[24][26] ), .QN(n368) );
  DFFRX1 \register_r_reg[24][25]  ( .D(n1892), .CK(clk), .RN(n3362), .Q(
        \register_r[24][25] ), .QN(n369) );
  DFFRX1 \register_r_reg[24][24]  ( .D(n1891), .CK(clk), .RN(n3362), .Q(
        \register_r[24][24] ), .QN(n370) );
  DFFRX1 \register_r_reg[24][23]  ( .D(n1890), .CK(clk), .RN(n3362), .Q(
        \register_r[24][23] ), .QN(n371) );
  DFFRX1 \register_r_reg[24][22]  ( .D(n1889), .CK(clk), .RN(n3362), .Q(
        \register_r[24][22] ), .QN(n372) );
  DFFRX1 \register_r_reg[24][21]  ( .D(n1888), .CK(clk), .RN(n3362), .Q(
        \register_r[24][21] ), .QN(n373) );
  DFFRX1 \register_r_reg[24][20]  ( .D(n1887), .CK(clk), .RN(n3362), .Q(
        \register_r[24][20] ), .QN(n374) );
  DFFRX1 \register_r_reg[24][19]  ( .D(n1886), .CK(clk), .RN(n3361), .Q(
        \register_r[24][19] ), .QN(n375) );
  DFFRX1 \register_r_reg[24][18]  ( .D(n1885), .CK(clk), .RN(n3361), .Q(
        \register_r[24][18] ), .QN(n376) );
  DFFRX1 \register_r_reg[24][17]  ( .D(n1884), .CK(clk), .RN(n3361), .Q(
        \register_r[24][17] ), .QN(n377) );
  DFFRX1 \register_r_reg[24][16]  ( .D(n1883), .CK(clk), .RN(n3361), .Q(
        \register_r[24][16] ), .QN(n378) );
  DFFRX1 \register_r_reg[24][15]  ( .D(n1882), .CK(clk), .RN(n3361), .Q(
        \register_r[24][15] ), .QN(n379) );
  DFFRX1 \register_r_reg[24][14]  ( .D(n1881), .CK(clk), .RN(n3361), .Q(
        \register_r[24][14] ), .QN(n380) );
  DFFRX1 \register_r_reg[24][13]  ( .D(n1880), .CK(clk), .RN(n3361), .Q(
        \register_r[24][13] ), .QN(n381) );
  DFFRX1 \register_r_reg[24][12]  ( .D(n1879), .CK(clk), .RN(n3361), .Q(
        \register_r[24][12] ), .QN(n382) );
  DFFRX1 \register_r_reg[24][11]  ( .D(n1878), .CK(clk), .RN(n3361), .Q(
        \register_r[24][11] ), .QN(n383) );
  DFFRX1 \register_r_reg[24][10]  ( .D(n1877), .CK(clk), .RN(n3361), .Q(
        \register_r[24][10] ), .QN(n384) );
  DFFRX1 \register_r_reg[24][9]  ( .D(n1876), .CK(clk), .RN(n3361), .Q(
        \register_r[24][9] ), .QN(n385) );
  DFFRX1 \register_r_reg[24][8]  ( .D(n1875), .CK(clk), .RN(n3361), .Q(
        \register_r[24][8] ), .QN(n386) );
  DFFRX1 \register_r_reg[24][7]  ( .D(n1874), .CK(clk), .RN(n3360), .Q(
        \register_r[24][7] ), .QN(n387) );
  DFFRX1 \register_r_reg[24][6]  ( .D(n1873), .CK(clk), .RN(n3360), .Q(
        \register_r[24][6] ), .QN(n388) );
  DFFRX1 \register_r_reg[24][5]  ( .D(n1872), .CK(clk), .RN(n3360), .Q(
        \register_r[24][5] ), .QN(n389) );
  DFFRX1 \register_r_reg[24][4]  ( .D(n1871), .CK(clk), .RN(n3360), .Q(
        \register_r[24][4] ), .QN(n390) );
  DFFRX1 \register_r_reg[24][3]  ( .D(n1870), .CK(clk), .RN(n3360), .Q(
        \register_r[24][3] ), .QN(n391) );
  DFFRX1 \register_r_reg[24][2]  ( .D(n1869), .CK(clk), .RN(n3360), .Q(
        \register_r[24][2] ), .QN(n392) );
  DFFRX1 \register_r_reg[24][1]  ( .D(n1868), .CK(clk), .RN(n3360), .Q(
        \register_r[24][1] ), .QN(n393) );
  DFFRX1 \register_r_reg[24][0]  ( .D(n1867), .CK(clk), .RN(n3360), .Q(
        \register_r[24][0] ), .QN(n394) );
  DFFRX1 \register_r_reg[20][23]  ( .D(n1762), .CK(clk), .RN(n3351), .Q(
        \register_r[20][23] ), .QN(n499) );
  DFFRX1 \register_r_reg[20][22]  ( .D(n1761), .CK(clk), .RN(n3351), .Q(
        \register_r[20][22] ), .QN(n500) );
  DFFRX1 \register_r_reg[20][21]  ( .D(n1760), .CK(clk), .RN(n3351), .Q(
        \register_r[20][21] ), .QN(n501) );
  DFFRX1 \register_r_reg[20][20]  ( .D(n1759), .CK(clk), .RN(n3351), .Q(
        \register_r[20][20] ), .QN(n502) );
  DFFRX1 \register_r_reg[20][19]  ( .D(n1758), .CK(clk), .RN(n3351), .Q(
        \register_r[20][19] ), .QN(n503) );
  DFFRX1 \register_r_reg[20][18]  ( .D(n1757), .CK(clk), .RN(n3351), .Q(
        \register_r[20][18] ), .QN(n504) );
  DFFRX1 \register_r_reg[20][17]  ( .D(n1756), .CK(clk), .RN(n3351), .Q(
        \register_r[20][17] ), .QN(n505) );
  DFFRX1 \register_r_reg[20][16]  ( .D(n1755), .CK(clk), .RN(n3351), .Q(
        \register_r[20][16] ), .QN(n506) );
  DFFRX1 \register_r_reg[20][15]  ( .D(n1754), .CK(clk), .RN(n3350), .Q(
        \register_r[20][15] ), .QN(n507) );
  DFFRX1 \register_r_reg[20][14]  ( .D(n1753), .CK(clk), .RN(n3350), .Q(
        \register_r[20][14] ), .QN(n508) );
  DFFRX1 \register_r_reg[20][13]  ( .D(n1752), .CK(clk), .RN(n3350), .Q(
        \register_r[20][13] ), .QN(n509) );
  DFFRX1 \register_r_reg[20][12]  ( .D(n1751), .CK(clk), .RN(n3350), .Q(
        \register_r[20][12] ), .QN(n510) );
  DFFRX1 \register_r_reg[20][11]  ( .D(n1750), .CK(clk), .RN(n3350), .Q(
        \register_r[20][11] ), .QN(n511) );
  DFFRX1 \register_r_reg[20][10]  ( .D(n1749), .CK(clk), .RN(n3350), .Q(
        \register_r[20][10] ), .QN(n512) );
  DFFRX1 \register_r_reg[20][9]  ( .D(n1748), .CK(clk), .RN(n3350), .Q(
        \register_r[20][9] ), .QN(n513) );
  DFFRX1 \register_r_reg[20][8]  ( .D(n1747), .CK(clk), .RN(n3350), .Q(
        \register_r[20][8] ), .QN(n514) );
  DFFRX1 \register_r_reg[20][7]  ( .D(n1746), .CK(clk), .RN(n3350), .Q(
        \register_r[20][7] ), .QN(n515) );
  DFFRX1 \register_r_reg[20][6]  ( .D(n1745), .CK(clk), .RN(n3350), .Q(
        \register_r[20][6] ), .QN(n516) );
  DFFRX1 \register_r_reg[20][5]  ( .D(n1744), .CK(clk), .RN(n3350), .Q(
        \register_r[20][5] ), .QN(n517) );
  DFFRX1 \register_r_reg[20][4]  ( .D(n1743), .CK(clk), .RN(n3350), .Q(
        \register_r[20][4] ), .QN(n518) );
  DFFRX1 \register_r_reg[20][3]  ( .D(n1742), .CK(clk), .RN(n3349), .Q(
        \register_r[20][3] ), .QN(n519) );
  DFFRX1 \register_r_reg[20][2]  ( .D(n1741), .CK(clk), .RN(n3349), .Q(
        \register_r[20][2] ), .QN(n520) );
  DFFRX1 \register_r_reg[20][1]  ( .D(n1740), .CK(clk), .RN(n3349), .Q(
        \register_r[20][1] ), .QN(n521) );
  DFFRX1 \register_r_reg[20][0]  ( .D(n1739), .CK(clk), .RN(n3349), .Q(
        \register_r[20][0] ), .QN(n522) );
  DFFRX1 \register_r_reg[16][23]  ( .D(n1634), .CK(clk), .RN(n3340), .Q(
        \register_r[16][23] ), .QN(n627) );
  DFFRX1 \register_r_reg[16][22]  ( .D(n1633), .CK(clk), .RN(n3340), .Q(
        \register_r[16][22] ), .QN(n628) );
  DFFRX1 \register_r_reg[16][21]  ( .D(n1632), .CK(clk), .RN(n3340), .Q(
        \register_r[16][21] ), .QN(n629) );
  DFFRX1 \register_r_reg[16][20]  ( .D(n1631), .CK(clk), .RN(n3340), .Q(
        \register_r[16][20] ), .QN(n630) );
  DFFRX1 \register_r_reg[16][19]  ( .D(n1630), .CK(clk), .RN(n3340), .Q(
        \register_r[16][19] ), .QN(n631) );
  DFFRX1 \register_r_reg[16][18]  ( .D(n1629), .CK(clk), .RN(n3340), .Q(
        \register_r[16][18] ), .QN(n632) );
  DFFRX1 \register_r_reg[16][17]  ( .D(n1628), .CK(clk), .RN(n3340), .Q(
        \register_r[16][17] ), .QN(n633) );
  DFFRX1 \register_r_reg[16][16]  ( .D(n1627), .CK(clk), .RN(n3340), .Q(
        \register_r[16][16] ), .QN(n634) );
  DFFRX1 \register_r_reg[16][15]  ( .D(n1626), .CK(clk), .RN(n3340), .Q(
        \register_r[16][15] ), .QN(n635) );
  DFFRX1 \register_r_reg[16][14]  ( .D(n1625), .CK(clk), .RN(n3340), .Q(
        \register_r[16][14] ), .QN(n636) );
  DFFRX1 \register_r_reg[16][13]  ( .D(n1624), .CK(clk), .RN(n3340), .Q(
        \register_r[16][13] ), .QN(n637) );
  DFFRX1 \register_r_reg[16][12]  ( .D(n1623), .CK(clk), .RN(n3340), .Q(
        \register_r[16][12] ), .QN(n638) );
  DFFRX1 \register_r_reg[16][11]  ( .D(n1622), .CK(clk), .RN(n3339), .Q(
        \register_r[16][11] ), .QN(n639) );
  DFFRX1 \register_r_reg[16][10]  ( .D(n1621), .CK(clk), .RN(n3339), .Q(
        \register_r[16][10] ), .QN(n640) );
  DFFRX1 \register_r_reg[16][9]  ( .D(n1620), .CK(clk), .RN(n3339), .Q(
        \register_r[16][9] ), .QN(n641) );
  DFFRX1 \register_r_reg[16][8]  ( .D(n1619), .CK(clk), .RN(n3339), .Q(
        \register_r[16][8] ), .QN(n642) );
  DFFRX1 \register_r_reg[16][7]  ( .D(n1618), .CK(clk), .RN(n3339), .Q(
        \register_r[16][7] ), .QN(n643) );
  DFFRX1 \register_r_reg[16][6]  ( .D(n1617), .CK(clk), .RN(n3339), .Q(
        \register_r[16][6] ), .QN(n644) );
  DFFRX1 \register_r_reg[16][5]  ( .D(n1616), .CK(clk), .RN(n3339), .Q(
        \register_r[16][5] ), .QN(n645) );
  DFFRX1 \register_r_reg[16][4]  ( .D(n1615), .CK(clk), .RN(n3339), .Q(
        \register_r[16][4] ), .QN(n646) );
  DFFRX1 \register_r_reg[16][3]  ( .D(n1614), .CK(clk), .RN(n3339), .Q(
        \register_r[16][3] ), .QN(n647) );
  DFFRX1 \register_r_reg[16][2]  ( .D(n1613), .CK(clk), .RN(n3339), .Q(
        \register_r[16][2] ), .QN(n648) );
  DFFRX1 \register_r_reg[16][1]  ( .D(n1612), .CK(clk), .RN(n3339), .Q(
        \register_r[16][1] ), .QN(n649) );
  DFFRX1 \register_r_reg[16][0]  ( .D(n1611), .CK(clk), .RN(n3339), .Q(
        \register_r[16][0] ), .QN(n650) );
  DFFRX1 \register_r_reg[12][31]  ( .D(n1514), .CK(clk), .RN(n3330), .Q(
        r_12[31]), .QN(n747) );
  DFFRX1 \register_r_reg[12][30]  ( .D(n1513), .CK(clk), .RN(n3330), .Q(
        r_12[30]), .QN(n748) );
  DFFRX1 \register_r_reg[12][29]  ( .D(n1512), .CK(clk), .RN(n3330), .Q(
        r_12[29]), .QN(n749) );
  DFFRX1 \register_r_reg[12][28]  ( .D(n1511), .CK(clk), .RN(n3330), .Q(
        r_12[28]), .QN(n750) );
  DFFRX1 \register_r_reg[12][27]  ( .D(n1510), .CK(clk), .RN(n3330), .Q(
        r_12[27]), .QN(n751) );
  DFFRX1 \register_r_reg[12][26]  ( .D(n1509), .CK(clk), .RN(n3330), .Q(
        r_12[26]), .QN(n752) );
  DFFRX1 \register_r_reg[12][25]  ( .D(n1508), .CK(clk), .RN(n3330), .Q(
        r_12[25]), .QN(n753) );
  DFFRX1 \register_r_reg[12][24]  ( .D(n1507), .CK(clk), .RN(n3330), .Q(
        r_12[24]), .QN(n754) );
  DFFRX1 \register_r_reg[12][23]  ( .D(n1506), .CK(clk), .RN(n3330), .Q(
        r_12[23]), .QN(n755) );
  DFFRX1 \register_r_reg[12][22]  ( .D(n1505), .CK(clk), .RN(n3330), .Q(
        r_12[22]), .QN(n756) );
  DFFRX1 \register_r_reg[12][21]  ( .D(n1504), .CK(clk), .RN(n3330), .Q(
        r_12[21]), .QN(n757) );
  DFFRX1 \register_r_reg[12][20]  ( .D(n1503), .CK(clk), .RN(n3330), .Q(
        r_12[20]), .QN(n758) );
  DFFRX1 \register_r_reg[12][19]  ( .D(n1502), .CK(clk), .RN(n3329), .Q(
        r_12[19]), .QN(n759) );
  DFFRX1 \register_r_reg[12][18]  ( .D(n1501), .CK(clk), .RN(n3329), .Q(
        r_12[18]), .QN(n760) );
  DFFRX1 \register_r_reg[12][17]  ( .D(n1500), .CK(clk), .RN(n3329), .Q(
        r_12[17]), .QN(n761) );
  DFFRX1 \register_r_reg[12][16]  ( .D(n1499), .CK(clk), .RN(n3329), .Q(
        r_12[16]), .QN(n762) );
  DFFRX1 \register_r_reg[12][15]  ( .D(n1498), .CK(clk), .RN(n3329), .Q(
        r_12[15]), .QN(n763) );
  DFFRX1 \register_r_reg[12][14]  ( .D(n1497), .CK(clk), .RN(n3329), .Q(
        r_12[14]), .QN(n764) );
  DFFRX1 \register_r_reg[12][13]  ( .D(n1496), .CK(clk), .RN(n3329), .Q(
        r_12[13]), .QN(n765) );
  DFFRX1 \register_r_reg[12][12]  ( .D(n1495), .CK(clk), .RN(n3329), .Q(
        r_12[12]), .QN(n766) );
  DFFRX1 \register_r_reg[12][11]  ( .D(n1494), .CK(clk), .RN(n3329), .Q(
        r_12[11]), .QN(n767) );
  DFFRX1 \register_r_reg[12][10]  ( .D(n1493), .CK(clk), .RN(n3329), .Q(
        r_12[10]), .QN(n768) );
  DFFRX1 \register_r_reg[12][9]  ( .D(n1492), .CK(clk), .RN(n3329), .Q(r_12[9]), .QN(n769) );
  DFFRX1 \register_r_reg[12][8]  ( .D(n1491), .CK(clk), .RN(n3329), .Q(r_12[8]), .QN(n770) );
  DFFRX1 \register_r_reg[12][7]  ( .D(n1490), .CK(clk), .RN(n3328), .Q(r_12[7]), .QN(n771) );
  DFFRX1 \register_r_reg[12][6]  ( .D(n1489), .CK(clk), .RN(n3328), .Q(r_12[6]), .QN(n772) );
  DFFRX1 \register_r_reg[12][5]  ( .D(n1488), .CK(clk), .RN(n3328), .Q(r_12[5]), .QN(n773) );
  DFFRX1 \register_r_reg[12][4]  ( .D(n1487), .CK(clk), .RN(n3328), .Q(r_12[4]), .QN(n774) );
  DFFRX1 \register_r_reg[12][3]  ( .D(n1486), .CK(clk), .RN(n3328), .Q(r_12[3]), .QN(n775) );
  DFFRX1 \register_r_reg[12][2]  ( .D(n1485), .CK(clk), .RN(n3328), .Q(r_12[2]), .QN(n776) );
  DFFRX1 \register_r_reg[12][1]  ( .D(n1484), .CK(clk), .RN(n3328), .Q(r_12[1]), .QN(n777) );
  DFFRX1 \register_r_reg[12][0]  ( .D(n1483), .CK(clk), .RN(n3328), .Q(r_12[0]), .QN(n778) );
  DFFRX1 \register_r_reg[8][31]  ( .D(n1386), .CK(clk), .RN(n3320), .Q(
        \register_r[8][31] ), .QN(n875) );
  DFFRX1 \register_r_reg[8][30]  ( .D(n1385), .CK(clk), .RN(n3320), .Q(
        \register_r[8][30] ), .QN(n876) );
  DFFRX1 \register_r_reg[8][29]  ( .D(n1384), .CK(clk), .RN(n3320), .Q(
        \register_r[8][29] ), .QN(n877) );
  DFFRX1 \register_r_reg[8][28]  ( .D(n1383), .CK(clk), .RN(n3320), .Q(
        \register_r[8][28] ), .QN(n878) );
  DFFRX1 \register_r_reg[8][27]  ( .D(n1382), .CK(clk), .RN(n3319), .Q(
        \register_r[8][27] ), .QN(n879) );
  DFFRX1 \register_r_reg[8][26]  ( .D(n1381), .CK(clk), .RN(n3319), .Q(
        \register_r[8][26] ), .QN(n880) );
  DFFRX1 \register_r_reg[8][25]  ( .D(n1380), .CK(clk), .RN(n3319), .Q(
        \register_r[8][25] ), .QN(n881) );
  DFFRX1 \register_r_reg[8][24]  ( .D(n1379), .CK(clk), .RN(n3319), .Q(
        \register_r[8][24] ), .QN(n882) );
  DFFRX1 \register_r_reg[8][23]  ( .D(n1378), .CK(clk), .RN(n3319), .Q(
        \register_r[8][23] ), .QN(n883) );
  DFFRX1 \register_r_reg[8][22]  ( .D(n1377), .CK(clk), .RN(n3319), .Q(
        \register_r[8][22] ), .QN(n884) );
  DFFRX1 \register_r_reg[8][21]  ( .D(n1376), .CK(clk), .RN(n3319), .Q(
        \register_r[8][21] ), .QN(n885) );
  DFFRX1 \register_r_reg[8][20]  ( .D(n1375), .CK(clk), .RN(n3319), .Q(
        \register_r[8][20] ), .QN(n886) );
  DFFRX1 \register_r_reg[8][19]  ( .D(n1374), .CK(clk), .RN(n3319), .Q(
        \register_r[8][19] ), .QN(n887) );
  DFFRX1 \register_r_reg[8][18]  ( .D(n1373), .CK(clk), .RN(n3319), .Q(
        \register_r[8][18] ), .QN(n888) );
  DFFRX1 \register_r_reg[8][17]  ( .D(n1372), .CK(clk), .RN(n3319), .Q(
        \register_r[8][17] ), .QN(n889) );
  DFFRX1 \register_r_reg[8][16]  ( .D(n1371), .CK(clk), .RN(n3319), .Q(
        \register_r[8][16] ), .QN(n890) );
  DFFRX1 \register_r_reg[8][15]  ( .D(n1370), .CK(clk), .RN(n3318), .Q(
        \register_r[8][15] ), .QN(n891) );
  DFFRX1 \register_r_reg[8][14]  ( .D(n1369), .CK(clk), .RN(n3318), .Q(
        \register_r[8][14] ), .QN(n892) );
  DFFRX1 \register_r_reg[8][13]  ( .D(n1368), .CK(clk), .RN(n3318), .Q(
        \register_r[8][13] ), .QN(n893) );
  DFFRX1 \register_r_reg[8][12]  ( .D(n1367), .CK(clk), .RN(n3318), .Q(
        \register_r[8][12] ), .QN(n894) );
  DFFRX1 \register_r_reg[8][11]  ( .D(n1366), .CK(clk), .RN(n3318), .Q(
        \register_r[8][11] ), .QN(n895) );
  DFFRX1 \register_r_reg[8][10]  ( .D(n1365), .CK(clk), .RN(n3318), .Q(
        \register_r[8][10] ), .QN(n896) );
  DFFRX1 \register_r_reg[8][9]  ( .D(n1364), .CK(clk), .RN(n3318), .Q(
        \register_r[8][9] ), .QN(n897) );
  DFFRX1 \register_r_reg[8][8]  ( .D(n1363), .CK(clk), .RN(n3318), .Q(
        \register_r[8][8] ), .QN(n898) );
  DFFRX1 \register_r_reg[8][7]  ( .D(n1362), .CK(clk), .RN(n3318), .Q(
        \register_r[8][7] ), .QN(n899) );
  DFFRX1 \register_r_reg[8][6]  ( .D(n1361), .CK(clk), .RN(n3318), .Q(
        \register_r[8][6] ), .QN(n900) );
  DFFRX1 \register_r_reg[8][5]  ( .D(n1360), .CK(clk), .RN(n3318), .Q(
        \register_r[8][5] ), .QN(n901) );
  DFFRX1 \register_r_reg[8][4]  ( .D(n1359), .CK(clk), .RN(n3318), .Q(
        \register_r[8][4] ), .QN(n902) );
  DFFRX1 \register_r_reg[8][3]  ( .D(n1358), .CK(clk), .RN(n3317), .Q(
        \register_r[8][3] ), .QN(n903) );
  DFFRX1 \register_r_reg[8][2]  ( .D(n1357), .CK(clk), .RN(n3317), .Q(
        \register_r[8][2] ), .QN(n904) );
  DFFRX1 \register_r_reg[8][1]  ( .D(n1356), .CK(clk), .RN(n3317), .Q(
        \register_r[8][1] ), .QN(n905) );
  DFFRX1 \register_r_reg[8][0]  ( .D(n1355), .CK(clk), .RN(n3317), .Q(
        \register_r[8][0] ), .QN(n906) );
  DFFRX1 \register_r_reg[4][31]  ( .D(n1258), .CK(clk), .RN(n3309), .Q(
        \register_r[4][31] ), .QN(n1003) );
  DFFRX1 \register_r_reg[4][30]  ( .D(n1257), .CK(clk), .RN(n3309), .Q(
        \register_r[4][30] ), .QN(n1004) );
  DFFRX1 \register_r_reg[4][29]  ( .D(n1256), .CK(clk), .RN(n3309), .Q(
        \register_r[4][29] ), .QN(n1005) );
  DFFRX1 \register_r_reg[4][28]  ( .D(n1255), .CK(clk), .RN(n3309), .Q(
        \register_r[4][28] ), .QN(n1006) );
  DFFRX1 \register_r_reg[4][27]  ( .D(n1254), .CK(clk), .RN(n3309), .Q(
        \register_r[4][27] ), .QN(n1007) );
  DFFRX1 \register_r_reg[4][26]  ( .D(n1253), .CK(clk), .RN(n3309), .Q(
        \register_r[4][26] ), .QN(n1008) );
  DFFRX1 \register_r_reg[4][25]  ( .D(n1252), .CK(clk), .RN(n3309), .Q(
        \register_r[4][25] ), .QN(n1009) );
  DFFRX1 \register_r_reg[4][24]  ( .D(n1251), .CK(clk), .RN(n3309), .Q(
        \register_r[4][24] ), .QN(n1010) );
  DFFRX1 \register_r_reg[4][23]  ( .D(n1250), .CK(clk), .RN(n3308), .Q(
        \register_r[4][23] ), .QN(n1011) );
  DFFRX1 \register_r_reg[4][22]  ( .D(n1249), .CK(clk), .RN(n3308), .Q(
        \register_r[4][22] ), .QN(n1012) );
  DFFRX1 \register_r_reg[4][21]  ( .D(n1248), .CK(clk), .RN(n3308), .Q(
        \register_r[4][21] ), .QN(n1013) );
  DFFRX1 \register_r_reg[4][20]  ( .D(n1247), .CK(clk), .RN(n3308), .Q(
        \register_r[4][20] ), .QN(n1014) );
  DFFRX1 \register_r_reg[4][19]  ( .D(n1246), .CK(clk), .RN(n3308), .Q(
        \register_r[4][19] ), .QN(n1015) );
  DFFRX1 \register_r_reg[4][18]  ( .D(n1245), .CK(clk), .RN(n3308), .Q(
        \register_r[4][18] ), .QN(n1016) );
  DFFRX1 \register_r_reg[4][17]  ( .D(n1244), .CK(clk), .RN(n3308), .Q(
        \register_r[4][17] ), .QN(n1017) );
  DFFRX1 \register_r_reg[4][16]  ( .D(n1243), .CK(clk), .RN(n3308), .Q(
        \register_r[4][16] ), .QN(n1018) );
  DFFRX1 \register_r_reg[4][15]  ( .D(n1242), .CK(clk), .RN(n3308), .Q(
        \register_r[4][15] ), .QN(n1019) );
  DFFRX1 \register_r_reg[4][14]  ( .D(n1241), .CK(clk), .RN(n3308), .Q(
        \register_r[4][14] ), .QN(n1020) );
  DFFRX1 \register_r_reg[4][13]  ( .D(n1240), .CK(clk), .RN(n3308), .Q(
        \register_r[4][13] ), .QN(n1021) );
  DFFRX1 \register_r_reg[4][12]  ( .D(n1239), .CK(clk), .RN(n3308), .Q(
        \register_r[4][12] ), .QN(n1022) );
  DFFRX1 \register_r_reg[4][11]  ( .D(n1238), .CK(clk), .RN(n3307), .Q(
        \register_r[4][11] ), .QN(n1023) );
  DFFRX1 \register_r_reg[4][10]  ( .D(n1237), .CK(clk), .RN(n3307), .Q(
        \register_r[4][10] ), .QN(n1024) );
  DFFRX1 \register_r_reg[4][9]  ( .D(n1236), .CK(clk), .RN(n3307), .Q(
        \register_r[4][9] ), .QN(n1025) );
  DFFRX1 \register_r_reg[4][8]  ( .D(n1235), .CK(clk), .RN(n3307), .Q(
        \register_r[4][8] ), .QN(n1026) );
  DFFRX1 \register_r_reg[4][7]  ( .D(n1234), .CK(clk), .RN(n3307), .Q(
        \register_r[4][7] ), .QN(n1027) );
  DFFRX1 \register_r_reg[4][6]  ( .D(n1233), .CK(clk), .RN(n3307), .Q(
        \register_r[4][6] ), .QN(n1028) );
  DFFRX1 \register_r_reg[4][5]  ( .D(n1232), .CK(clk), .RN(n3307), .Q(
        \register_r[4][5] ), .QN(n1029) );
  DFFRX1 \register_r_reg[4][4]  ( .D(n1231), .CK(clk), .RN(n3307), .Q(
        \register_r[4][4] ), .QN(n1030) );
  DFFRX1 \register_r_reg[4][3]  ( .D(n1230), .CK(clk), .RN(n3307), .Q(
        \register_r[4][3] ), .QN(n1031) );
  DFFRX1 \register_r_reg[4][2]  ( .D(n1229), .CK(clk), .RN(n3307), .Q(
        \register_r[4][2] ), .QN(n1032) );
  DFFRX1 \register_r_reg[4][1]  ( .D(n1228), .CK(clk), .RN(n3307), .Q(
        \register_r[4][1] ), .QN(n1033) );
  DFFRX1 \register_r_reg[4][0]  ( .D(n1227), .CK(clk), .RN(n3307), .Q(
        \register_r[4][0] ), .QN(n1034) );
  DFFRX1 \register_r_reg[30][31]  ( .D(n2090), .CK(clk), .RN(n3378), .Q(
        \register_r[30][31] ), .QN(n171) );
  DFFRX1 \register_r_reg[30][30]  ( .D(n2089), .CK(clk), .RN(n3378), .Q(
        \register_r[30][30] ), .QN(n172) );
  DFFRX1 \register_r_reg[30][29]  ( .D(n2088), .CK(clk), .RN(n3378), .Q(
        \register_r[30][29] ), .QN(n173) );
  DFFRX1 \register_r_reg[30][28]  ( .D(n2087), .CK(clk), .RN(n3378), .Q(
        \register_r[30][28] ), .QN(n174) );
  DFFRX1 \register_r_reg[30][27]  ( .D(n2086), .CK(clk), .RN(n3378), .Q(
        \register_r[30][27] ), .QN(n175) );
  DFFRX1 \register_r_reg[30][26]  ( .D(n2085), .CK(clk), .RN(n3378), .Q(
        \register_r[30][26] ), .QN(n176) );
  DFFRX1 \register_r_reg[30][25]  ( .D(n2084), .CK(clk), .RN(n3378), .Q(
        \register_r[30][25] ), .QN(n177) );
  DFFRX1 \register_r_reg[30][24]  ( .D(n2083), .CK(clk), .RN(n3378), .Q(
        \register_r[30][24] ), .QN(n178) );
  DFFRX1 \register_r_reg[30][23]  ( .D(n2082), .CK(clk), .RN(n3378), .Q(
        \register_r[30][23] ), .QN(n179) );
  DFFRX1 \register_r_reg[30][22]  ( .D(n2081), .CK(clk), .RN(n3378), .Q(
        \register_r[30][22] ), .QN(n180) );
  DFFRX1 \register_r_reg[30][21]  ( .D(n2080), .CK(clk), .RN(n3378), .Q(
        \register_r[30][21] ), .QN(n181) );
  DFFRX1 \register_r_reg[30][20]  ( .D(n2079), .CK(clk), .RN(n3378), .Q(
        \register_r[30][20] ), .QN(n182) );
  DFFRX1 \register_r_reg[30][19]  ( .D(n2078), .CK(clk), .RN(n3377), .Q(
        \register_r[30][19] ), .QN(n183) );
  DFFRX1 \register_r_reg[30][18]  ( .D(n2077), .CK(clk), .RN(n3377), .Q(
        \register_r[30][18] ), .QN(n184) );
  DFFRX1 \register_r_reg[30][17]  ( .D(n2076), .CK(clk), .RN(n3377), .Q(
        \register_r[30][17] ), .QN(n185) );
  DFFRX1 \register_r_reg[30][16]  ( .D(n2075), .CK(clk), .RN(n3377), .Q(
        \register_r[30][16] ), .QN(n186) );
  DFFRX1 \register_r_reg[30][15]  ( .D(n2074), .CK(clk), .RN(n3377), .Q(
        \register_r[30][15] ), .QN(n187) );
  DFFRX1 \register_r_reg[30][14]  ( .D(n2073), .CK(clk), .RN(n3377), .Q(
        \register_r[30][14] ), .QN(n188) );
  DFFRX1 \register_r_reg[30][13]  ( .D(n2072), .CK(clk), .RN(n3377), .Q(
        \register_r[30][13] ), .QN(n189) );
  DFFRX1 \register_r_reg[30][12]  ( .D(n2071), .CK(clk), .RN(n3377), .Q(
        \register_r[30][12] ), .QN(n190) );
  DFFRX1 \register_r_reg[30][11]  ( .D(n2070), .CK(clk), .RN(n3377), .Q(
        \register_r[30][11] ), .QN(n191) );
  DFFRX1 \register_r_reg[30][10]  ( .D(n2069), .CK(clk), .RN(n3377), .Q(
        \register_r[30][10] ), .QN(n192) );
  DFFRX1 \register_r_reg[30][9]  ( .D(n2068), .CK(clk), .RN(n3377), .Q(
        \register_r[30][9] ), .QN(n193) );
  DFFRX1 \register_r_reg[30][8]  ( .D(n2067), .CK(clk), .RN(n3377), .Q(
        \register_r[30][8] ), .QN(n194) );
  DFFRX1 \register_r_reg[30][7]  ( .D(n2066), .CK(clk), .RN(n3376), .Q(
        \register_r[30][7] ), .QN(n195) );
  DFFRX1 \register_r_reg[30][6]  ( .D(n2065), .CK(clk), .RN(n3376), .Q(
        \register_r[30][6] ), .QN(n196) );
  DFFRX1 \register_r_reg[30][5]  ( .D(n2064), .CK(clk), .RN(n3376), .Q(
        \register_r[30][5] ), .QN(n197) );
  DFFRX1 \register_r_reg[30][4]  ( .D(n2063), .CK(clk), .RN(n3376), .Q(
        \register_r[30][4] ), .QN(n198) );
  DFFRX1 \register_r_reg[30][3]  ( .D(n2062), .CK(clk), .RN(n3376), .Q(
        \register_r[30][3] ), .QN(n199) );
  DFFRX1 \register_r_reg[30][2]  ( .D(n2061), .CK(clk), .RN(n3376), .Q(
        \register_r[30][2] ), .QN(n200) );
  DFFRX1 \register_r_reg[30][1]  ( .D(n2060), .CK(clk), .RN(n3376), .Q(
        \register_r[30][1] ), .QN(n201) );
  DFFRX1 \register_r_reg[30][0]  ( .D(n2059), .CK(clk), .RN(n3376), .Q(
        \register_r[30][0] ), .QN(n202) );
  DFFRX1 \register_r_reg[26][31]  ( .D(n1962), .CK(clk), .RN(n3368), .Q(
        \register_r[26][31] ), .QN(n299) );
  DFFRX1 \register_r_reg[26][30]  ( .D(n1961), .CK(clk), .RN(n3368), .Q(
        \register_r[26][30] ), .QN(n300) );
  DFFRX1 \register_r_reg[26][29]  ( .D(n1960), .CK(clk), .RN(n3368), .Q(
        \register_r[26][29] ), .QN(n301) );
  DFFRX1 \register_r_reg[26][28]  ( .D(n1959), .CK(clk), .RN(n3368), .Q(
        \register_r[26][28] ), .QN(n302) );
  DFFRX1 \register_r_reg[26][27]  ( .D(n1958), .CK(clk), .RN(n3367), .Q(
        \register_r[26][27] ), .QN(n303) );
  DFFRX1 \register_r_reg[26][26]  ( .D(n1957), .CK(clk), .RN(n3367), .Q(
        \register_r[26][26] ), .QN(n304) );
  DFFRX1 \register_r_reg[26][25]  ( .D(n1956), .CK(clk), .RN(n3367), .Q(
        \register_r[26][25] ), .QN(n305) );
  DFFRX1 \register_r_reg[26][24]  ( .D(n1955), .CK(clk), .RN(n3367), .Q(
        \register_r[26][24] ), .QN(n306) );
  DFFRX1 \register_r_reg[26][23]  ( .D(n1954), .CK(clk), .RN(n3367), .Q(
        \register_r[26][23] ), .QN(n307) );
  DFFRX1 \register_r_reg[26][22]  ( .D(n1953), .CK(clk), .RN(n3367), .Q(
        \register_r[26][22] ), .QN(n308) );
  DFFRX1 \register_r_reg[26][21]  ( .D(n1952), .CK(clk), .RN(n3367), .Q(
        \register_r[26][21] ), .QN(n309) );
  DFFRX1 \register_r_reg[26][20]  ( .D(n1951), .CK(clk), .RN(n3367), .Q(
        \register_r[26][20] ), .QN(n310) );
  DFFRX1 \register_r_reg[26][19]  ( .D(n1950), .CK(clk), .RN(n3367), .Q(
        \register_r[26][19] ), .QN(n311) );
  DFFRX1 \register_r_reg[26][18]  ( .D(n1949), .CK(clk), .RN(n3367), .Q(
        \register_r[26][18] ), .QN(n312) );
  DFFRX1 \register_r_reg[26][17]  ( .D(n1948), .CK(clk), .RN(n3367), .Q(
        \register_r[26][17] ), .QN(n313) );
  DFFRX1 \register_r_reg[26][16]  ( .D(n1947), .CK(clk), .RN(n3367), .Q(
        \register_r[26][16] ), .QN(n314) );
  DFFRX1 \register_r_reg[26][15]  ( .D(n1946), .CK(clk), .RN(n3366), .Q(
        \register_r[26][15] ), .QN(n315) );
  DFFRX1 \register_r_reg[26][14]  ( .D(n1945), .CK(clk), .RN(n3366), .Q(
        \register_r[26][14] ), .QN(n316) );
  DFFRX1 \register_r_reg[26][13]  ( .D(n1944), .CK(clk), .RN(n3366), .Q(
        \register_r[26][13] ), .QN(n317) );
  DFFRX1 \register_r_reg[26][12]  ( .D(n1943), .CK(clk), .RN(n3366), .Q(
        \register_r[26][12] ), .QN(n318) );
  DFFRX1 \register_r_reg[26][11]  ( .D(n1942), .CK(clk), .RN(n3366), .Q(
        \register_r[26][11] ), .QN(n319) );
  DFFRX1 \register_r_reg[26][10]  ( .D(n1941), .CK(clk), .RN(n3366), .Q(
        \register_r[26][10] ), .QN(n320) );
  DFFRX1 \register_r_reg[26][9]  ( .D(n1940), .CK(clk), .RN(n3366), .Q(
        \register_r[26][9] ), .QN(n321) );
  DFFRX1 \register_r_reg[26][8]  ( .D(n1939), .CK(clk), .RN(n3366), .Q(
        \register_r[26][8] ), .QN(n322) );
  DFFRX1 \register_r_reg[26][7]  ( .D(n1938), .CK(clk), .RN(n3366), .Q(
        \register_r[26][7] ), .QN(n323) );
  DFFRX1 \register_r_reg[26][6]  ( .D(n1937), .CK(clk), .RN(n3366), .Q(
        \register_r[26][6] ), .QN(n324) );
  DFFRX1 \register_r_reg[26][5]  ( .D(n1936), .CK(clk), .RN(n3366), .Q(
        \register_r[26][5] ), .QN(n325) );
  DFFRX1 \register_r_reg[26][4]  ( .D(n1935), .CK(clk), .RN(n3366), .Q(
        \register_r[26][4] ), .QN(n326) );
  DFFRX1 \register_r_reg[26][3]  ( .D(n1934), .CK(clk), .RN(n3365), .Q(
        \register_r[26][3] ), .QN(n327) );
  DFFRX1 \register_r_reg[26][2]  ( .D(n1933), .CK(clk), .RN(n3365), .Q(
        \register_r[26][2] ), .QN(n328) );
  DFFRX1 \register_r_reg[26][1]  ( .D(n1932), .CK(clk), .RN(n3365), .Q(
        \register_r[26][1] ), .QN(n329) );
  DFFRX1 \register_r_reg[26][0]  ( .D(n1931), .CK(clk), .RN(n3365), .Q(
        \register_r[26][0] ), .QN(n330) );
  DFFRX1 \register_r_reg[22][23]  ( .D(n1826), .CK(clk), .RN(n3356), .Q(
        \register_r[22][23] ), .QN(n435) );
  DFFRX1 \register_r_reg[22][22]  ( .D(n1825), .CK(clk), .RN(n3356), .Q(
        \register_r[22][22] ), .QN(n436) );
  DFFRX1 \register_r_reg[22][21]  ( .D(n1824), .CK(clk), .RN(n3356), .Q(
        \register_r[22][21] ), .QN(n437) );
  DFFRX1 \register_r_reg[22][20]  ( .D(n1823), .CK(clk), .RN(n3356), .Q(
        \register_r[22][20] ), .QN(n438) );
  DFFRX1 \register_r_reg[22][19]  ( .D(n1822), .CK(clk), .RN(n3356), .Q(
        \register_r[22][19] ), .QN(n439) );
  DFFRX1 \register_r_reg[22][18]  ( .D(n1821), .CK(clk), .RN(n3356), .Q(
        \register_r[22][18] ), .QN(n440) );
  DFFRX1 \register_r_reg[22][17]  ( .D(n1820), .CK(clk), .RN(n3356), .Q(
        \register_r[22][17] ), .QN(n441) );
  DFFRX1 \register_r_reg[22][16]  ( .D(n1819), .CK(clk), .RN(n3356), .Q(
        \register_r[22][16] ), .QN(n442) );
  DFFRX1 \register_r_reg[22][15]  ( .D(n1818), .CK(clk), .RN(n3356), .Q(
        \register_r[22][15] ), .QN(n443) );
  DFFRX1 \register_r_reg[22][14]  ( .D(n1817), .CK(clk), .RN(n3356), .Q(
        \register_r[22][14] ), .QN(n444) );
  DFFRX1 \register_r_reg[22][13]  ( .D(n1816), .CK(clk), .RN(n3356), .Q(
        \register_r[22][13] ), .QN(n445) );
  DFFRX1 \register_r_reg[22][12]  ( .D(n1815), .CK(clk), .RN(n3356), .Q(
        \register_r[22][12] ), .QN(n446) );
  DFFRX1 \register_r_reg[22][11]  ( .D(n1814), .CK(clk), .RN(n3355), .Q(
        \register_r[22][11] ), .QN(n447) );
  DFFRX1 \register_r_reg[22][10]  ( .D(n1813), .CK(clk), .RN(n3355), .Q(
        \register_r[22][10] ), .QN(n448) );
  DFFRX1 \register_r_reg[22][9]  ( .D(n1812), .CK(clk), .RN(n3355), .Q(
        \register_r[22][9] ), .QN(n449) );
  DFFRX1 \register_r_reg[22][8]  ( .D(n1811), .CK(clk), .RN(n3355), .Q(
        \register_r[22][8] ), .QN(n450) );
  DFFRX1 \register_r_reg[22][7]  ( .D(n1810), .CK(clk), .RN(n3355), .Q(
        \register_r[22][7] ), .QN(n451) );
  DFFRX1 \register_r_reg[22][6]  ( .D(n1809), .CK(clk), .RN(n3355), .Q(
        \register_r[22][6] ), .QN(n452) );
  DFFRX1 \register_r_reg[22][5]  ( .D(n1808), .CK(clk), .RN(n3355), .Q(
        \register_r[22][5] ), .QN(n453) );
  DFFRX1 \register_r_reg[22][4]  ( .D(n1807), .CK(clk), .RN(n3355), .Q(
        \register_r[22][4] ), .QN(n454) );
  DFFRX1 \register_r_reg[22][3]  ( .D(n1806), .CK(clk), .RN(n3355), .Q(
        \register_r[22][3] ), .QN(n455) );
  DFFRX1 \register_r_reg[22][2]  ( .D(n1805), .CK(clk), .RN(n3355), .Q(
        \register_r[22][2] ), .QN(n456) );
  DFFRX1 \register_r_reg[22][1]  ( .D(n1804), .CK(clk), .RN(n3355), .Q(
        \register_r[22][1] ), .QN(n457) );
  DFFRX1 \register_r_reg[22][0]  ( .D(n1803), .CK(clk), .RN(n3355), .Q(
        \register_r[22][0] ), .QN(n458) );
  DFFRX1 \register_r_reg[18][23]  ( .D(n1698), .CK(clk), .RN(n3346), .Q(
        \register_r[18][23] ), .QN(n563) );
  DFFRX1 \register_r_reg[18][22]  ( .D(n1697), .CK(clk), .RN(n3346), .Q(
        \register_r[18][22] ), .QN(n564) );
  DFFRX1 \register_r_reg[18][21]  ( .D(n1696), .CK(clk), .RN(n3346), .Q(
        \register_r[18][21] ), .QN(n565) );
  DFFRX1 \register_r_reg[18][20]  ( .D(n1695), .CK(clk), .RN(n3346), .Q(
        \register_r[18][20] ), .QN(n566) );
  DFFRX1 \register_r_reg[18][19]  ( .D(n1694), .CK(clk), .RN(n3345), .Q(
        \register_r[18][19] ), .QN(n567) );
  DFFRX1 \register_r_reg[18][18]  ( .D(n1693), .CK(clk), .RN(n3345), .Q(
        \register_r[18][18] ), .QN(n568) );
  DFFRX1 \register_r_reg[18][17]  ( .D(n1692), .CK(clk), .RN(n3345), .Q(
        \register_r[18][17] ), .QN(n569) );
  DFFRX1 \register_r_reg[18][16]  ( .D(n1691), .CK(clk), .RN(n3345), .Q(
        \register_r[18][16] ), .QN(n570) );
  DFFRX1 \register_r_reg[18][15]  ( .D(n1690), .CK(clk), .RN(n3345), .Q(
        \register_r[18][15] ), .QN(n571) );
  DFFRX1 \register_r_reg[18][14]  ( .D(n1689), .CK(clk), .RN(n3345), .Q(
        \register_r[18][14] ), .QN(n572) );
  DFFRX1 \register_r_reg[18][13]  ( .D(n1688), .CK(clk), .RN(n3345), .Q(
        \register_r[18][13] ), .QN(n573) );
  DFFRX1 \register_r_reg[18][12]  ( .D(n1687), .CK(clk), .RN(n3345), .Q(
        \register_r[18][12] ), .QN(n574) );
  DFFRX1 \register_r_reg[18][11]  ( .D(n1686), .CK(clk), .RN(n3345), .Q(
        \register_r[18][11] ), .QN(n575) );
  DFFRX1 \register_r_reg[18][10]  ( .D(n1685), .CK(clk), .RN(n3345), .Q(
        \register_r[18][10] ), .QN(n576) );
  DFFRX1 \register_r_reg[18][9]  ( .D(n1684), .CK(clk), .RN(n3345), .Q(
        \register_r[18][9] ), .QN(n577) );
  DFFRX1 \register_r_reg[18][8]  ( .D(n1683), .CK(clk), .RN(n3345), .Q(
        \register_r[18][8] ), .QN(n578) );
  DFFRX1 \register_r_reg[18][7]  ( .D(n1682), .CK(clk), .RN(n3344), .Q(
        \register_r[18][7] ), .QN(n579) );
  DFFRX1 \register_r_reg[18][6]  ( .D(n1681), .CK(clk), .RN(n3344), .Q(
        \register_r[18][6] ), .QN(n580) );
  DFFRX1 \register_r_reg[18][5]  ( .D(n1680), .CK(clk), .RN(n3344), .Q(
        \register_r[18][5] ), .QN(n581) );
  DFFRX1 \register_r_reg[18][4]  ( .D(n1679), .CK(clk), .RN(n3344), .Q(
        \register_r[18][4] ), .QN(n582) );
  DFFRX1 \register_r_reg[18][3]  ( .D(n1678), .CK(clk), .RN(n3344), .Q(
        \register_r[18][3] ), .QN(n583) );
  DFFRX1 \register_r_reg[18][2]  ( .D(n1677), .CK(clk), .RN(n3344), .Q(
        \register_r[18][2] ), .QN(n584) );
  DFFRX1 \register_r_reg[18][1]  ( .D(n1676), .CK(clk), .RN(n3344), .Q(
        \register_r[18][1] ), .QN(n585) );
  DFFRX1 \register_r_reg[18][0]  ( .D(n1675), .CK(clk), .RN(n3344), .Q(
        \register_r[18][0] ), .QN(n586) );
  DFFRX1 \register_r_reg[14][31]  ( .D(n1578), .CK(clk), .RN(n3336), .Q(
        \register_r[14][31] ), .QN(n683) );
  DFFRX1 \register_r_reg[14][30]  ( .D(n1577), .CK(clk), .RN(n3336), .Q(
        \register_r[14][30] ), .QN(n684) );
  DFFRX1 \register_r_reg[14][29]  ( .D(n1576), .CK(clk), .RN(n3336), .Q(
        \register_r[14][29] ), .QN(n685) );
  DFFRX1 \register_r_reg[14][28]  ( .D(n1575), .CK(clk), .RN(n3336), .Q(
        \register_r[14][28] ), .QN(n686) );
  DFFRX1 \register_r_reg[14][27]  ( .D(n1574), .CK(clk), .RN(n3335), .Q(
        \register_r[14][27] ), .QN(n687) );
  DFFRX1 \register_r_reg[14][26]  ( .D(n1573), .CK(clk), .RN(n3335), .Q(
        \register_r[14][26] ), .QN(n688) );
  DFFRX1 \register_r_reg[14][25]  ( .D(n1572), .CK(clk), .RN(n3335), .Q(
        \register_r[14][25] ), .QN(n689) );
  DFFRX1 \register_r_reg[14][24]  ( .D(n1571), .CK(clk), .RN(n3335), .Q(
        \register_r[14][24] ), .QN(n690) );
  DFFRX1 \register_r_reg[14][23]  ( .D(n1570), .CK(clk), .RN(n3335), .Q(
        \register_r[14][23] ), .QN(n691) );
  DFFRX1 \register_r_reg[14][22]  ( .D(n1569), .CK(clk), .RN(n3335), .Q(
        \register_r[14][22] ), .QN(n692) );
  DFFRX1 \register_r_reg[14][21]  ( .D(n1568), .CK(clk), .RN(n3335), .Q(
        \register_r[14][21] ), .QN(n693) );
  DFFRX1 \register_r_reg[14][20]  ( .D(n1567), .CK(clk), .RN(n3335), .Q(
        \register_r[14][20] ), .QN(n694) );
  DFFRX1 \register_r_reg[14][19]  ( .D(n1566), .CK(clk), .RN(n3335), .Q(
        \register_r[14][19] ), .QN(n695) );
  DFFRX1 \register_r_reg[14][18]  ( .D(n1565), .CK(clk), .RN(n3335), .Q(
        \register_r[14][18] ), .QN(n696) );
  DFFRX1 \register_r_reg[14][17]  ( .D(n1564), .CK(clk), .RN(n3335), .Q(
        \register_r[14][17] ), .QN(n697) );
  DFFRX1 \register_r_reg[14][16]  ( .D(n1563), .CK(clk), .RN(n3335), .Q(
        \register_r[14][16] ), .QN(n698) );
  DFFRX1 \register_r_reg[14][15]  ( .D(n1562), .CK(clk), .RN(n3334), .Q(
        \register_r[14][15] ), .QN(n699) );
  DFFRX1 \register_r_reg[14][14]  ( .D(n1561), .CK(clk), .RN(n3334), .Q(
        \register_r[14][14] ), .QN(n700) );
  DFFRX1 \register_r_reg[14][13]  ( .D(n1560), .CK(clk), .RN(n3334), .Q(
        \register_r[14][13] ), .QN(n701) );
  DFFRX1 \register_r_reg[14][12]  ( .D(n1559), .CK(clk), .RN(n3334), .Q(
        \register_r[14][12] ), .QN(n702) );
  DFFRX1 \register_r_reg[14][11]  ( .D(n1558), .CK(clk), .RN(n3334), .Q(
        \register_r[14][11] ), .QN(n703) );
  DFFRX1 \register_r_reg[14][10]  ( .D(n1557), .CK(clk), .RN(n3334), .Q(
        \register_r[14][10] ), .QN(n704) );
  DFFRX1 \register_r_reg[14][9]  ( .D(n1556), .CK(clk), .RN(n3334), .Q(
        \register_r[14][9] ), .QN(n705) );
  DFFRX1 \register_r_reg[14][8]  ( .D(n1555), .CK(clk), .RN(n3334), .Q(
        \register_r[14][8] ), .QN(n706) );
  DFFRX1 \register_r_reg[14][7]  ( .D(n1554), .CK(clk), .RN(n3334), .Q(
        \register_r[14][7] ), .QN(n707) );
  DFFRX1 \register_r_reg[14][6]  ( .D(n1553), .CK(clk), .RN(n3334), .Q(
        \register_r[14][6] ), .QN(n708) );
  DFFRX1 \register_r_reg[14][5]  ( .D(n1552), .CK(clk), .RN(n3334), .Q(
        \register_r[14][5] ), .QN(n709) );
  DFFRX1 \register_r_reg[14][4]  ( .D(n1551), .CK(clk), .RN(n3334), .Q(
        \register_r[14][4] ), .QN(n710) );
  DFFRX1 \register_r_reg[14][3]  ( .D(n1550), .CK(clk), .RN(n3333), .Q(
        \register_r[14][3] ), .QN(n711) );
  DFFRX1 \register_r_reg[14][2]  ( .D(n1549), .CK(clk), .RN(n3333), .Q(
        \register_r[14][2] ), .QN(n712) );
  DFFRX1 \register_r_reg[14][1]  ( .D(n1548), .CK(clk), .RN(n3333), .Q(
        \register_r[14][1] ), .QN(n713) );
  DFFRX1 \register_r_reg[14][0]  ( .D(n1547), .CK(clk), .RN(n3333), .Q(
        \register_r[14][0] ), .QN(n714) );
  DFFRX1 \register_r_reg[10][31]  ( .D(n1450), .CK(clk), .RN(n3325), .Q(
        \register_r[10][31] ), .QN(n811) );
  DFFRX1 \register_r_reg[10][30]  ( .D(n1449), .CK(clk), .RN(n3325), .Q(
        \register_r[10][30] ), .QN(n812) );
  DFFRX1 \register_r_reg[10][29]  ( .D(n1448), .CK(clk), .RN(n3325), .Q(
        \register_r[10][29] ), .QN(n813) );
  DFFRX1 \register_r_reg[10][28]  ( .D(n1447), .CK(clk), .RN(n3325), .Q(
        \register_r[10][28] ), .QN(n814) );
  DFFRX1 \register_r_reg[10][27]  ( .D(n1446), .CK(clk), .RN(n3325), .Q(
        \register_r[10][27] ), .QN(n815) );
  DFFRX1 \register_r_reg[10][26]  ( .D(n1445), .CK(clk), .RN(n3325), .Q(
        \register_r[10][26] ), .QN(n816) );
  DFFRX1 \register_r_reg[10][25]  ( .D(n1444), .CK(clk), .RN(n3325), .Q(
        \register_r[10][25] ), .QN(n817) );
  DFFRX1 \register_r_reg[10][24]  ( .D(n1443), .CK(clk), .RN(n3325), .Q(
        \register_r[10][24] ), .QN(n818) );
  DFFRX1 \register_r_reg[10][23]  ( .D(n1442), .CK(clk), .RN(n3324), .Q(
        \register_r[10][23] ), .QN(n819) );
  DFFRX1 \register_r_reg[10][22]  ( .D(n1441), .CK(clk), .RN(n3324), .Q(
        \register_r[10][22] ), .QN(n820) );
  DFFRX1 \register_r_reg[10][21]  ( .D(n1440), .CK(clk), .RN(n3324), .Q(
        \register_r[10][21] ), .QN(n821) );
  DFFRX1 \register_r_reg[10][20]  ( .D(n1439), .CK(clk), .RN(n3324), .Q(
        \register_r[10][20] ), .QN(n822) );
  DFFRX1 \register_r_reg[10][19]  ( .D(n1438), .CK(clk), .RN(n3324), .Q(
        \register_r[10][19] ), .QN(n823) );
  DFFRX1 \register_r_reg[10][18]  ( .D(n1437), .CK(clk), .RN(n3324), .Q(
        \register_r[10][18] ), .QN(n824) );
  DFFRX1 \register_r_reg[10][17]  ( .D(n1436), .CK(clk), .RN(n3324), .Q(
        \register_r[10][17] ), .QN(n825) );
  DFFRX1 \register_r_reg[10][16]  ( .D(n1435), .CK(clk), .RN(n3324), .Q(
        \register_r[10][16] ), .QN(n826) );
  DFFRX1 \register_r_reg[10][15]  ( .D(n1434), .CK(clk), .RN(n3324), .Q(
        \register_r[10][15] ), .QN(n827) );
  DFFRX1 \register_r_reg[10][14]  ( .D(n1433), .CK(clk), .RN(n3324), .Q(
        \register_r[10][14] ), .QN(n828) );
  DFFRX1 \register_r_reg[10][13]  ( .D(n1432), .CK(clk), .RN(n3324), .Q(
        \register_r[10][13] ), .QN(n829) );
  DFFRX1 \register_r_reg[10][12]  ( .D(n1431), .CK(clk), .RN(n3324), .Q(
        \register_r[10][12] ), .QN(n830) );
  DFFRX1 \register_r_reg[10][11]  ( .D(n1430), .CK(clk), .RN(n3323), .Q(
        \register_r[10][11] ), .QN(n831) );
  DFFRX1 \register_r_reg[10][10]  ( .D(n1429), .CK(clk), .RN(n3323), .Q(
        \register_r[10][10] ), .QN(n832) );
  DFFRX1 \register_r_reg[10][9]  ( .D(n1428), .CK(clk), .RN(n3323), .Q(
        \register_r[10][9] ), .QN(n833) );
  DFFRX1 \register_r_reg[10][8]  ( .D(n1427), .CK(clk), .RN(n3323), .Q(
        \register_r[10][8] ), .QN(n834) );
  DFFRX1 \register_r_reg[10][7]  ( .D(n1426), .CK(clk), .RN(n3323), .Q(
        \register_r[10][7] ), .QN(n835) );
  DFFRX1 \register_r_reg[10][6]  ( .D(n1425), .CK(clk), .RN(n3323), .Q(
        \register_r[10][6] ), .QN(n836) );
  DFFRX1 \register_r_reg[10][5]  ( .D(n1424), .CK(clk), .RN(n3323), .Q(
        \register_r[10][5] ), .QN(n837) );
  DFFRX1 \register_r_reg[10][4]  ( .D(n1423), .CK(clk), .RN(n3323), .Q(
        \register_r[10][4] ), .QN(n838) );
  DFFRX1 \register_r_reg[10][3]  ( .D(n1422), .CK(clk), .RN(n3323), .Q(
        \register_r[10][3] ), .QN(n839) );
  DFFRX1 \register_r_reg[10][2]  ( .D(n1421), .CK(clk), .RN(n3323), .Q(
        \register_r[10][2] ), .QN(n840) );
  DFFRX1 \register_r_reg[10][1]  ( .D(n1420), .CK(clk), .RN(n3323), .Q(
        \register_r[10][1] ), .QN(n841) );
  DFFRX1 \register_r_reg[10][0]  ( .D(n1419), .CK(clk), .RN(n3323), .Q(
        \register_r[10][0] ), .QN(n842) );
  DFFRX1 \register_r_reg[6][31]  ( .D(n1322), .CK(clk), .RN(n3314), .Q(
        \register_r[6][31] ), .QN(n939) );
  DFFRX1 \register_r_reg[6][30]  ( .D(n1321), .CK(clk), .RN(n3314), .Q(
        \register_r[6][30] ), .QN(n940) );
  DFFRX1 \register_r_reg[6][29]  ( .D(n1320), .CK(clk), .RN(n3314), .Q(
        \register_r[6][29] ), .QN(n941) );
  DFFRX1 \register_r_reg[6][28]  ( .D(n1319), .CK(clk), .RN(n3314), .Q(
        \register_r[6][28] ), .QN(n942) );
  DFFRX1 \register_r_reg[6][27]  ( .D(n1318), .CK(clk), .RN(n3314), .Q(
        \register_r[6][27] ), .QN(n943) );
  DFFRX1 \register_r_reg[6][26]  ( .D(n1317), .CK(clk), .RN(n3314), .Q(
        \register_r[6][26] ), .QN(n944) );
  DFFRX1 \register_r_reg[6][25]  ( .D(n1316), .CK(clk), .RN(n3314), .Q(
        \register_r[6][25] ), .QN(n945) );
  DFFRX1 \register_r_reg[6][24]  ( .D(n1315), .CK(clk), .RN(n3314), .Q(
        \register_r[6][24] ), .QN(n946) );
  DFFRX1 \register_r_reg[6][23]  ( .D(n1314), .CK(clk), .RN(n3314), .Q(
        \register_r[6][23] ), .QN(n947) );
  DFFRX1 \register_r_reg[6][22]  ( .D(n1313), .CK(clk), .RN(n3314), .Q(
        \register_r[6][22] ), .QN(n948) );
  DFFRX1 \register_r_reg[6][21]  ( .D(n1312), .CK(clk), .RN(n3314), .Q(
        \register_r[6][21] ), .QN(n949) );
  DFFRX1 \register_r_reg[6][20]  ( .D(n1311), .CK(clk), .RN(n3314), .Q(
        \register_r[6][20] ), .QN(n950) );
  DFFRX1 \register_r_reg[6][19]  ( .D(n1310), .CK(clk), .RN(n3313), .Q(
        \register_r[6][19] ), .QN(n951) );
  DFFRX1 \register_r_reg[6][18]  ( .D(n1309), .CK(clk), .RN(n3313), .Q(
        \register_r[6][18] ), .QN(n952) );
  DFFRX1 \register_r_reg[6][17]  ( .D(n1308), .CK(clk), .RN(n3313), .Q(
        \register_r[6][17] ), .QN(n953) );
  DFFRX1 \register_r_reg[6][16]  ( .D(n1307), .CK(clk), .RN(n3313), .Q(
        \register_r[6][16] ), .QN(n954) );
  DFFRX1 \register_r_reg[6][15]  ( .D(n1306), .CK(clk), .RN(n3313), .Q(
        \register_r[6][15] ), .QN(n955) );
  DFFRX1 \register_r_reg[6][14]  ( .D(n1305), .CK(clk), .RN(n3313), .Q(
        \register_r[6][14] ), .QN(n956) );
  DFFRX1 \register_r_reg[6][13]  ( .D(n1304), .CK(clk), .RN(n3313), .Q(
        \register_r[6][13] ), .QN(n957) );
  DFFRX1 \register_r_reg[6][12]  ( .D(n1303), .CK(clk), .RN(n3313), .Q(
        \register_r[6][12] ), .QN(n958) );
  DFFRX1 \register_r_reg[6][11]  ( .D(n1302), .CK(clk), .RN(n3313), .Q(
        \register_r[6][11] ), .QN(n959) );
  DFFRX1 \register_r_reg[6][10]  ( .D(n1301), .CK(clk), .RN(n3313), .Q(
        \register_r[6][10] ), .QN(n960) );
  DFFRX1 \register_r_reg[6][9]  ( .D(n1300), .CK(clk), .RN(n3313), .Q(
        \register_r[6][9] ), .QN(n961) );
  DFFRX1 \register_r_reg[6][8]  ( .D(n1299), .CK(clk), .RN(n3313), .Q(
        \register_r[6][8] ), .QN(n962) );
  DFFRX1 \register_r_reg[6][7]  ( .D(n1298), .CK(clk), .RN(n3312), .Q(
        \register_r[6][7] ), .QN(n963) );
  DFFRX1 \register_r_reg[6][6]  ( .D(n1297), .CK(clk), .RN(n3312), .Q(
        \register_r[6][6] ), .QN(n964) );
  DFFRX1 \register_r_reg[6][5]  ( .D(n1296), .CK(clk), .RN(n3312), .Q(
        \register_r[6][5] ), .QN(n965) );
  DFFRX1 \register_r_reg[6][4]  ( .D(n1295), .CK(clk), .RN(n3312), .Q(
        \register_r[6][4] ), .QN(n966) );
  DFFRX1 \register_r_reg[6][3]  ( .D(n1294), .CK(clk), .RN(n3312), .Q(
        \register_r[6][3] ), .QN(n967) );
  DFFRX1 \register_r_reg[6][2]  ( .D(n1293), .CK(clk), .RN(n3312), .Q(
        \register_r[6][2] ), .QN(n968) );
  DFFRX1 \register_r_reg[6][1]  ( .D(n1292), .CK(clk), .RN(n3312), .Q(
        \register_r[6][1] ), .QN(n969) );
  DFFRX1 \register_r_reg[6][0]  ( .D(n1291), .CK(clk), .RN(n3312), .Q(
        \register_r[6][0] ), .QN(n970) );
  DFFRX1 \register_r_reg[3][31]  ( .D(n1226), .CK(clk), .RN(n3306), .Q(
        \register_r[3][31] ), .QN(n1035) );
  DFFRX1 \register_r_reg[3][30]  ( .D(n1225), .CK(clk), .RN(n3306), .Q(
        \register_r[3][30] ), .QN(n1036) );
  DFFRX1 \register_r_reg[3][29]  ( .D(n1224), .CK(clk), .RN(n3306), .Q(
        \register_r[3][29] ), .QN(n1037) );
  DFFRX1 \register_r_reg[3][28]  ( .D(n1223), .CK(clk), .RN(n3306), .Q(
        \register_r[3][28] ), .QN(n1038) );
  DFFRX1 \register_r_reg[3][27]  ( .D(n1222), .CK(clk), .RN(n3306), .Q(
        \register_r[3][27] ), .QN(n1039) );
  DFFRX1 \register_r_reg[3][26]  ( .D(n1221), .CK(clk), .RN(n3306), .Q(
        \register_r[3][26] ), .QN(n1040) );
  DFFRX1 \register_r_reg[3][25]  ( .D(n1220), .CK(clk), .RN(n3306), .Q(
        \register_r[3][25] ), .QN(n1041) );
  DFFRX1 \register_r_reg[3][24]  ( .D(n1219), .CK(clk), .RN(n3306), .Q(
        \register_r[3][24] ), .QN(n1042) );
  DFFRX1 \register_r_reg[3][23]  ( .D(n1218), .CK(clk), .RN(n3306), .Q(
        \register_r[3][23] ), .QN(n1043) );
  DFFRX1 \register_r_reg[3][22]  ( .D(n1217), .CK(clk), .RN(n3306), .Q(
        \register_r[3][22] ), .QN(n1044) );
  DFFRX1 \register_r_reg[3][21]  ( .D(n1216), .CK(clk), .RN(n3306), .Q(
        \register_r[3][21] ), .QN(n1045) );
  DFFRX1 \register_r_reg[3][20]  ( .D(n1215), .CK(clk), .RN(n3306), .Q(
        \register_r[3][20] ), .QN(n1046) );
  DFFRX1 \register_r_reg[3][19]  ( .D(n1214), .CK(clk), .RN(n3305), .Q(
        \register_r[3][19] ), .QN(n1047) );
  DFFRX1 \register_r_reg[3][18]  ( .D(n1213), .CK(clk), .RN(n3305), .Q(
        \register_r[3][18] ), .QN(n1048) );
  DFFRX1 \register_r_reg[3][17]  ( .D(n1212), .CK(clk), .RN(n3305), .Q(
        \register_r[3][17] ), .QN(n1049) );
  DFFRX1 \register_r_reg[3][16]  ( .D(n1211), .CK(clk), .RN(n3305), .Q(
        \register_r[3][16] ), .QN(n1050) );
  DFFRX1 \register_r_reg[3][15]  ( .D(n1210), .CK(clk), .RN(n3305), .Q(
        \register_r[3][15] ), .QN(n1051) );
  DFFRX1 \register_r_reg[3][14]  ( .D(n1209), .CK(clk), .RN(n3305), .Q(
        \register_r[3][14] ), .QN(n1052) );
  DFFRX1 \register_r_reg[3][13]  ( .D(n1208), .CK(clk), .RN(n3305), .Q(
        \register_r[3][13] ), .QN(n1053) );
  DFFRX1 \register_r_reg[3][12]  ( .D(n1207), .CK(clk), .RN(n3305), .Q(
        \register_r[3][12] ), .QN(n1054) );
  DFFRX1 \register_r_reg[3][11]  ( .D(n1206), .CK(clk), .RN(n3305), .Q(
        \register_r[3][11] ), .QN(n1055) );
  DFFRX1 \register_r_reg[3][10]  ( .D(n1205), .CK(clk), .RN(n3305), .Q(
        \register_r[3][10] ), .QN(n1056) );
  DFFRX1 \register_r_reg[3][9]  ( .D(n1204), .CK(clk), .RN(n3305), .Q(
        \register_r[3][9] ), .QN(n1057) );
  DFFRX1 \register_r_reg[3][8]  ( .D(n1203), .CK(clk), .RN(n3305), .Q(
        \register_r[3][8] ), .QN(n1058) );
  DFFRX1 \register_r_reg[3][7]  ( .D(n1202), .CK(clk), .RN(n3304), .Q(
        \register_r[3][7] ), .QN(n1059) );
  DFFRX1 \register_r_reg[3][6]  ( .D(n1201), .CK(clk), .RN(n3304), .Q(
        \register_r[3][6] ), .QN(n1060) );
  DFFRX1 \register_r_reg[3][5]  ( .D(n1200), .CK(clk), .RN(n3304), .Q(
        \register_r[3][5] ), .QN(n1061) );
  DFFRX1 \register_r_reg[3][4]  ( .D(n1199), .CK(clk), .RN(n3304), .Q(
        \register_r[3][4] ), .QN(n1062) );
  DFFRX1 \register_r_reg[3][3]  ( .D(n1198), .CK(clk), .RN(n3304), .Q(
        \register_r[3][3] ), .QN(n1063) );
  DFFRX1 \register_r_reg[3][2]  ( .D(n1197), .CK(clk), .RN(n3304), .Q(
        \register_r[3][2] ), .QN(n1064) );
  DFFRX1 \register_r_reg[3][1]  ( .D(n1196), .CK(clk), .RN(n3304), .Q(
        \register_r[3][1] ), .QN(n1065) );
  DFFRX1 \register_r_reg[3][0]  ( .D(n1195), .CK(clk), .RN(n3304), .Q(
        \register_r[3][0] ), .QN(n1066) );
  DFFRX1 \register_r_reg[1][31]  ( .D(n1162), .CK(clk), .RN(n3301), .Q(
        \register_r[1][31] ), .QN(n1099) );
  DFFRX1 \register_r_reg[1][30]  ( .D(n1161), .CK(clk), .RN(n3301), .Q(
        \register_r[1][30] ), .QN(n1100) );
  DFFRX1 \register_r_reg[1][29]  ( .D(n1160), .CK(clk), .RN(n3301), .Q(
        \register_r[1][29] ), .QN(n1101) );
  DFFRX1 \register_r_reg[1][28]  ( .D(n1159), .CK(clk), .RN(n3301), .Q(
        \register_r[1][28] ), .QN(n1102) );
  DFFRX1 \register_r_reg[1][27]  ( .D(n1158), .CK(clk), .RN(n3301), .Q(
        \register_r[1][27] ), .QN(n1103) );
  DFFRX1 \register_r_reg[1][26]  ( .D(n1157), .CK(clk), .RN(n3301), .Q(
        \register_r[1][26] ), .QN(n1104) );
  DFFRX1 \register_r_reg[1][25]  ( .D(n1156), .CK(clk), .RN(n3301), .Q(
        \register_r[1][25] ), .QN(n1105) );
  DFFRX1 \register_r_reg[1][24]  ( .D(n1155), .CK(clk), .RN(n3301), .Q(
        \register_r[1][24] ), .QN(n1106) );
  DFFRX1 \register_r_reg[1][23]  ( .D(n1154), .CK(clk), .RN(n3300), .Q(
        \register_r[1][23] ), .QN(n1107) );
  DFFRX1 \register_r_reg[1][22]  ( .D(n1153), .CK(clk), .RN(n3300), .Q(
        \register_r[1][22] ), .QN(n1108) );
  DFFRX1 \register_r_reg[1][21]  ( .D(n1152), .CK(clk), .RN(n3300), .Q(
        \register_r[1][21] ), .QN(n1109) );
  DFFRX1 \register_r_reg[1][20]  ( .D(n1151), .CK(clk), .RN(n3300), .Q(
        \register_r[1][20] ), .QN(n1110) );
  DFFRX1 \register_r_reg[1][19]  ( .D(n1150), .CK(clk), .RN(n3300), .Q(
        \register_r[1][19] ), .QN(n1111) );
  DFFRX1 \register_r_reg[1][18]  ( .D(n1149), .CK(clk), .RN(n3300), .Q(
        \register_r[1][18] ), .QN(n1112) );
  DFFRX1 \register_r_reg[1][17]  ( .D(n1148), .CK(clk), .RN(n3300), .Q(
        \register_r[1][17] ), .QN(n1113) );
  DFFRX1 \register_r_reg[1][16]  ( .D(n1147), .CK(clk), .RN(n3300), .Q(
        \register_r[1][16] ), .QN(n1114) );
  DFFRX1 \register_r_reg[1][15]  ( .D(n1146), .CK(clk), .RN(n3300), .Q(
        \register_r[1][15] ), .QN(n1115) );
  DFFRX1 \register_r_reg[1][14]  ( .D(n1145), .CK(clk), .RN(n3300), .Q(
        \register_r[1][14] ), .QN(n1116) );
  DFFRX1 \register_r_reg[1][13]  ( .D(n1144), .CK(clk), .RN(n3300), .Q(
        \register_r[1][13] ), .QN(n1117) );
  DFFRX1 \register_r_reg[1][12]  ( .D(n1143), .CK(clk), .RN(n3300), .Q(
        \register_r[1][12] ), .QN(n1118) );
  DFFRX1 \register_r_reg[1][11]  ( .D(n1142), .CK(clk), .RN(n3299), .Q(
        \register_r[1][11] ), .QN(n1119) );
  DFFRX1 \register_r_reg[1][10]  ( .D(n1141), .CK(clk), .RN(n3299), .Q(
        \register_r[1][10] ), .QN(n1120) );
  DFFRX1 \register_r_reg[1][9]  ( .D(n1140), .CK(clk), .RN(n3299), .Q(
        \register_r[1][9] ), .QN(n1121) );
  DFFRX1 \register_r_reg[1][8]  ( .D(n1139), .CK(clk), .RN(n3299), .Q(
        \register_r[1][8] ), .QN(n1122) );
  DFFRX1 \register_r_reg[1][7]  ( .D(n1138), .CK(clk), .RN(n3299), .Q(
        \register_r[1][7] ), .QN(n1123) );
  DFFRX1 \register_r_reg[1][6]  ( .D(n1137), .CK(clk), .RN(n3299), .Q(
        \register_r[1][6] ), .QN(n1124) );
  DFFRX1 \register_r_reg[1][5]  ( .D(n1136), .CK(clk), .RN(n3299), .Q(
        \register_r[1][5] ), .QN(n1125) );
  DFFRX1 \register_r_reg[1][4]  ( .D(n1135), .CK(clk), .RN(n3299), .Q(
        \register_r[1][4] ), .QN(n1126) );
  DFFRX1 \register_r_reg[1][3]  ( .D(n1134), .CK(clk), .RN(n3299), .Q(
        \register_r[1][3] ), .QN(n1127) );
  DFFRX1 \register_r_reg[1][2]  ( .D(n1133), .CK(clk), .RN(n3299), .Q(
        \register_r[1][2] ), .QN(n1128) );
  DFFRX1 \register_r_reg[1][1]  ( .D(n1132), .CK(clk), .RN(n3299), .Q(
        \register_r[1][1] ), .QN(n1129) );
  DFFRX1 \register_r_reg[1][0]  ( .D(n1131), .CK(clk), .RN(n3299), .Q(
        \register_r[1][0] ), .QN(n1130) );
  DFFRX1 \register_r_reg[22][31]  ( .D(n1834), .CK(clk), .RN(n3357), .Q(
        \register_r[22][31] ), .QN(n427) );
  DFFRX1 \register_r_reg[22][30]  ( .D(n1833), .CK(clk), .RN(n3357), .Q(
        \register_r[22][30] ), .QN(n428) );
  DFFRX1 \register_r_reg[22][29]  ( .D(n1832), .CK(clk), .RN(n3357), .Q(
        \register_r[22][29] ), .QN(n429) );
  DFFRX1 \register_r_reg[22][28]  ( .D(n1831), .CK(clk), .RN(n3357), .Q(
        \register_r[22][28] ), .QN(n430) );
  DFFRX1 \register_r_reg[22][27]  ( .D(n1830), .CK(clk), .RN(n3357), .Q(
        \register_r[22][27] ), .QN(n431) );
  DFFRX1 \register_r_reg[22][26]  ( .D(n1829), .CK(clk), .RN(n3357), .Q(
        \register_r[22][26] ), .QN(n432) );
  DFFRX1 \register_r_reg[22][25]  ( .D(n1828), .CK(clk), .RN(n3357), .Q(
        \register_r[22][25] ), .QN(n433) );
  DFFRX1 \register_r_reg[22][24]  ( .D(n1827), .CK(clk), .RN(n3357), .Q(
        \register_r[22][24] ), .QN(n434) );
  DFFRX1 \register_r_reg[23][31]  ( .D(n1866), .CK(clk), .RN(n3360), .Q(
        \register_r[23][31] ), .QN(n395) );
  DFFRX1 \register_r_reg[23][30]  ( .D(n1865), .CK(clk), .RN(n3360), .Q(
        \register_r[23][30] ), .QN(n396) );
  DFFRX1 \register_r_reg[23][29]  ( .D(n1864), .CK(clk), .RN(n3360), .Q(
        \register_r[23][29] ), .QN(n397) );
  DFFRX1 \register_r_reg[23][28]  ( .D(n1863), .CK(clk), .RN(n3360), .Q(
        \register_r[23][28] ), .QN(n398) );
  DFFRX1 \register_r_reg[23][27]  ( .D(n1862), .CK(clk), .RN(n3359), .Q(
        \register_r[23][27] ), .QN(n399) );
  DFFRX1 \register_r_reg[23][26]  ( .D(n1861), .CK(clk), .RN(n3359), .Q(
        \register_r[23][26] ), .QN(n400) );
  DFFRX1 \register_r_reg[23][25]  ( .D(n1860), .CK(clk), .RN(n3359), .Q(
        \register_r[23][25] ), .QN(n401) );
  DFFRX1 \register_r_reg[23][24]  ( .D(n1859), .CK(clk), .RN(n3359), .Q(
        \register_r[23][24] ), .QN(n402) );
  DFFRX1 \register_r_reg[21][31]  ( .D(n1802), .CK(clk), .RN(n3354), .Q(
        \register_r[21][31] ), .QN(n459) );
  DFFRX1 \register_r_reg[21][30]  ( .D(n1801), .CK(clk), .RN(n3354), .Q(
        \register_r[21][30] ), .QN(n460) );
  DFFRX1 \register_r_reg[21][29]  ( .D(n1800), .CK(clk), .RN(n3354), .Q(
        \register_r[21][29] ), .QN(n461) );
  DFFRX1 \register_r_reg[21][28]  ( .D(n1799), .CK(clk), .RN(n3354), .Q(
        \register_r[21][28] ), .QN(n462) );
  DFFRX1 \register_r_reg[21][27]  ( .D(n1798), .CK(clk), .RN(n3354), .Q(
        \register_r[21][27] ), .QN(n463) );
  DFFRX1 \register_r_reg[21][26]  ( .D(n1797), .CK(clk), .RN(n3354), .Q(
        \register_r[21][26] ), .QN(n464) );
  DFFRX1 \register_r_reg[21][25]  ( .D(n1796), .CK(clk), .RN(n3354), .Q(
        \register_r[21][25] ), .QN(n465) );
  DFFRX1 \register_r_reg[21][24]  ( .D(n1795), .CK(clk), .RN(n3354), .Q(
        \register_r[21][24] ), .QN(n466) );
  DFFRX1 \register_r_reg[20][31]  ( .D(n1770), .CK(clk), .RN(n3352), .Q(
        \register_r[20][31] ), .QN(n491) );
  DFFRX1 \register_r_reg[20][30]  ( .D(n1769), .CK(clk), .RN(n3352), .Q(
        \register_r[20][30] ), .QN(n492) );
  DFFRX1 \register_r_reg[20][29]  ( .D(n1768), .CK(clk), .RN(n3352), .Q(
        \register_r[20][29] ), .QN(n493) );
  DFFRX1 \register_r_reg[20][28]  ( .D(n1767), .CK(clk), .RN(n3352), .Q(
        \register_r[20][28] ), .QN(n494) );
  DFFRX1 \register_r_reg[20][27]  ( .D(n1766), .CK(clk), .RN(n3351), .Q(
        \register_r[20][27] ), .QN(n495) );
  DFFRX1 \register_r_reg[20][26]  ( .D(n1765), .CK(clk), .RN(n3351), .Q(
        \register_r[20][26] ), .QN(n496) );
  DFFRX1 \register_r_reg[20][25]  ( .D(n1764), .CK(clk), .RN(n3351), .Q(
        \register_r[20][25] ), .QN(n497) );
  DFFRX1 \register_r_reg[20][24]  ( .D(n1763), .CK(clk), .RN(n3351), .Q(
        \register_r[20][24] ), .QN(n498) );
  DFFRX1 \register_r_reg[18][31]  ( .D(n1706), .CK(clk), .RN(n3346), .Q(
        \register_r[18][31] ), .QN(n555) );
  DFFRX1 \register_r_reg[18][30]  ( .D(n1705), .CK(clk), .RN(n3346), .Q(
        \register_r[18][30] ), .QN(n556) );
  DFFRX1 \register_r_reg[18][29]  ( .D(n1704), .CK(clk), .RN(n3346), .Q(
        \register_r[18][29] ), .QN(n557) );
  DFFRX1 \register_r_reg[18][28]  ( .D(n1703), .CK(clk), .RN(n3346), .Q(
        \register_r[18][28] ), .QN(n558) );
  DFFRX1 \register_r_reg[18][27]  ( .D(n1702), .CK(clk), .RN(n3346), .Q(
        \register_r[18][27] ), .QN(n559) );
  DFFRX1 \register_r_reg[18][26]  ( .D(n1701), .CK(clk), .RN(n3346), .Q(
        \register_r[18][26] ), .QN(n560) );
  DFFRX1 \register_r_reg[18][25]  ( .D(n1700), .CK(clk), .RN(n3346), .Q(
        \register_r[18][25] ), .QN(n561) );
  DFFRX1 \register_r_reg[18][24]  ( .D(n1699), .CK(clk), .RN(n3346), .Q(
        \register_r[18][24] ), .QN(n562) );
  DFFRX1 \register_r_reg[16][31]  ( .D(n1642), .CK(clk), .RN(n3341), .Q(
        \register_r[16][31] ), .QN(n619) );
  DFFRX1 \register_r_reg[16][30]  ( .D(n1641), .CK(clk), .RN(n3341), .Q(
        \register_r[16][30] ), .QN(n620) );
  DFFRX1 \register_r_reg[16][29]  ( .D(n1640), .CK(clk), .RN(n3341), .Q(
        \register_r[16][29] ), .QN(n621) );
  DFFRX1 \register_r_reg[16][28]  ( .D(n1639), .CK(clk), .RN(n3341), .Q(
        \register_r[16][28] ), .QN(n622) );
  DFFRX1 \register_r_reg[16][27]  ( .D(n1638), .CK(clk), .RN(n3341), .Q(
        \register_r[16][27] ), .QN(n623) );
  DFFRX1 \register_r_reg[16][26]  ( .D(n1637), .CK(clk), .RN(n3341), .Q(
        \register_r[16][26] ), .QN(n624) );
  DFFRX1 \register_r_reg[16][25]  ( .D(n1636), .CK(clk), .RN(n3341), .Q(
        \register_r[16][25] ), .QN(n625) );
  DFFRX1 \register_r_reg[16][24]  ( .D(n1635), .CK(clk), .RN(n3341), .Q(
        \register_r[16][24] ), .QN(n626) );
  DFFRX1 \register_r_reg[19][31]  ( .D(n1738), .CK(clk), .RN(n3349), .Q(
        \register_r[19][31] ), .QN(n523) );
  DFFRX1 \register_r_reg[19][30]  ( .D(n1737), .CK(clk), .RN(n3349), .Q(
        \register_r[19][30] ), .QN(n524) );
  DFFRX1 \register_r_reg[19][29]  ( .D(n1736), .CK(clk), .RN(n3349), .Q(
        \register_r[19][29] ), .QN(n525) );
  DFFRX1 \register_r_reg[19][28]  ( .D(n1735), .CK(clk), .RN(n3349), .Q(
        \register_r[19][28] ), .QN(n526) );
  DFFRX1 \register_r_reg[19][27]  ( .D(n1734), .CK(clk), .RN(n3349), .Q(
        \register_r[19][27] ), .QN(n527) );
  DFFRX1 \register_r_reg[19][26]  ( .D(n1733), .CK(clk), .RN(n3349), .Q(
        \register_r[19][26] ), .QN(n528) );
  DFFRX1 \register_r_reg[19][25]  ( .D(n1732), .CK(clk), .RN(n3349), .Q(
        \register_r[19][25] ), .QN(n529) );
  DFFRX1 \register_r_reg[19][24]  ( .D(n1731), .CK(clk), .RN(n3349), .Q(
        \register_r[19][24] ), .QN(n530) );
  DFFRX1 \register_r_reg[17][31]  ( .D(n1674), .CK(clk), .RN(n3344), .Q(
        \register_r[17][31] ), .QN(n587) );
  DFFRX1 \register_r_reg[17][30]  ( .D(n1673), .CK(clk), .RN(n3344), .Q(
        \register_r[17][30] ), .QN(n588) );
  DFFRX1 \register_r_reg[17][29]  ( .D(n1672), .CK(clk), .RN(n3344), .Q(
        \register_r[17][29] ), .QN(n589) );
  DFFRX1 \register_r_reg[2][31]  ( .D(n1194), .CK(clk), .RN(n3304), .QN(n1067)
         );
  DFFRX1 \register_r_reg[2][30]  ( .D(n1193), .CK(clk), .RN(n3304), .QN(n1068)
         );
  DFFRX1 \register_r_reg[2][29]  ( .D(n1192), .CK(clk), .RN(n3304), .QN(n1069)
         );
  DFFRX1 \register_r_reg[2][28]  ( .D(n1191), .CK(clk), .RN(n3304), .QN(n1070)
         );
  DFFRX1 \register_r_reg[2][27]  ( .D(n1190), .CK(clk), .RN(n3303), .QN(n1071)
         );
  DFFRX1 \register_r_reg[2][26]  ( .D(n1189), .CK(clk), .RN(n3303), .QN(n1072)
         );
  DFFRX1 \register_r_reg[2][25]  ( .D(n1188), .CK(clk), .RN(n3303), .QN(n1073)
         );
  DFFRX1 \register_r_reg[2][24]  ( .D(n1187), .CK(clk), .RN(n3303), .QN(n1074)
         );
  DFFRX1 \register_r_reg[2][23]  ( .D(n1186), .CK(clk), .RN(n3303), .QN(n1075)
         );
  DFFRX1 \register_r_reg[2][22]  ( .D(n1185), .CK(clk), .RN(n3303), .QN(n1076)
         );
  DFFRX1 \register_r_reg[2][21]  ( .D(n1184), .CK(clk), .RN(n3303), .QN(n1077)
         );
  DFFRX1 \register_r_reg[2][20]  ( .D(n1183), .CK(clk), .RN(n3303), .QN(n1078)
         );
  DFFRX1 \register_r_reg[2][19]  ( .D(n1182), .CK(clk), .RN(n3303), .QN(n1079)
         );
  DFFRX1 \register_r_reg[2][18]  ( .D(n1181), .CK(clk), .RN(n3303), .QN(n1080)
         );
  DFFRX1 \register_r_reg[2][17]  ( .D(n1180), .CK(clk), .RN(n3303), .QN(n1081)
         );
  DFFRX1 \register_r_reg[2][16]  ( .D(n1179), .CK(clk), .RN(n3303), .QN(n1082)
         );
  DFFRX1 \register_r_reg[2][15]  ( .D(n1178), .CK(clk), .RN(n3302), .QN(n1083)
         );
  DFFRX1 \register_r_reg[2][14]  ( .D(n1177), .CK(clk), .RN(n3302), .QN(n1084)
         );
  DFFRX1 \register_r_reg[2][13]  ( .D(n1176), .CK(clk), .RN(n3302), .QN(n1085)
         );
  DFFRX1 \register_r_reg[2][12]  ( .D(n1175), .CK(clk), .RN(n3302), .QN(n1086)
         );
  DFFRX1 \register_r_reg[2][11]  ( .D(n1174), .CK(clk), .RN(n3302), .QN(n1087)
         );
  DFFRX1 \register_r_reg[2][10]  ( .D(n1173), .CK(clk), .RN(n3302), .QN(n1088)
         );
  DFFRX1 \register_r_reg[2][9]  ( .D(n1172), .CK(clk), .RN(n3302), .QN(n1089)
         );
  DFFRX1 \register_r_reg[2][8]  ( .D(n1171), .CK(clk), .RN(n3302), .QN(n1090)
         );
  DFFRX1 \register_r_reg[2][7]  ( .D(n1170), .CK(clk), .RN(n3302), .QN(n1091)
         );
  DFFRX1 \register_r_reg[2][6]  ( .D(n1169), .CK(clk), .RN(n3302), .QN(n1092)
         );
  DFFRX1 \register_r_reg[2][5]  ( .D(n1168), .CK(clk), .RN(n3302), .QN(n1093)
         );
  DFFRX1 \register_r_reg[2][4]  ( .D(n1167), .CK(clk), .RN(n3302), .QN(n1094)
         );
  DFFRX1 \register_r_reg[2][3]  ( .D(n1166), .CK(clk), .RN(n3301), .QN(n1095)
         );
  DFFRX1 \register_r_reg[2][2]  ( .D(n1165), .CK(clk), .RN(n3301), .QN(n1096)
         );
  DFFRX1 \register_r_reg[2][1]  ( .D(n1164), .CK(clk), .RN(n3301), .QN(n1097)
         );
  DFFRX1 \register_r_reg[2][0]  ( .D(n1163), .CK(clk), .RN(n3301), .QN(n1098)
         );
  CLKBUFX3 U3 ( .A(n3082), .Y(n3099) );
  CLKBUFX3 U4 ( .A(n2552), .Y(n2571) );
  CLKBUFX3 U5 ( .A(n3081), .Y(n3101) );
  CLKBUFX3 U6 ( .A(n3081), .Y(n3100) );
  CLKBUFX3 U7 ( .A(n2552), .Y(n2572) );
  CLKBUFX3 U8 ( .A(n2553), .Y(n2573) );
  CLKINVX1 U9 ( .A(WriteData[3]), .Y(n3436) );
  CLKINVX1 U10 ( .A(WriteData[4]), .Y(n3435) );
  CLKINVX1 U11 ( .A(WriteData[5]), .Y(n3434) );
  CLKINVX1 U12 ( .A(WriteData[6]), .Y(n3433) );
  CLKINVX1 U13 ( .A(WriteData[7]), .Y(n3432) );
  CLKINVX1 U14 ( .A(WriteData[8]), .Y(n3431) );
  CLKINVX1 U15 ( .A(WriteData[9]), .Y(n3430) );
  CLKINVX1 U16 ( .A(WriteData[31]), .Y(n3408) );
  CLKINVX1 U17 ( .A(WriteData[0]), .Y(n3439) );
  CLKINVX1 U18 ( .A(WriteData[1]), .Y(n3438) );
  CLKINVX1 U19 ( .A(WriteData[2]), .Y(n3437) );
  CLKINVX1 U20 ( .A(WriteData[10]), .Y(n3429) );
  CLKINVX1 U21 ( .A(WriteData[11]), .Y(n3428) );
  CLKINVX1 U22 ( .A(WriteData[12]), .Y(n3427) );
  CLKINVX1 U23 ( .A(WriteData[13]), .Y(n3426) );
  CLKINVX1 U24 ( .A(WriteData[14]), .Y(n3425) );
  CLKINVX1 U25 ( .A(WriteData[15]), .Y(n3424) );
  CLKINVX1 U26 ( .A(WriteData[16]), .Y(n3423) );
  CLKINVX1 U27 ( .A(WriteData[17]), .Y(n3422) );
  CLKINVX1 U28 ( .A(WriteData[18]), .Y(n3421) );
  CLKINVX1 U29 ( .A(WriteData[19]), .Y(n3420) );
  CLKINVX1 U30 ( .A(WriteData[20]), .Y(n3419) );
  CLKINVX1 U31 ( .A(WriteData[21]), .Y(n3418) );
  CLKINVX1 U32 ( .A(WriteData[22]), .Y(n3417) );
  CLKINVX1 U33 ( .A(WriteData[23]), .Y(n3416) );
  CLKINVX1 U34 ( .A(WriteData[24]), .Y(n3415) );
  CLKINVX1 U35 ( .A(WriteData[25]), .Y(n3414) );
  CLKINVX1 U36 ( .A(WriteData[26]), .Y(n3413) );
  CLKINVX1 U37 ( .A(WriteData[27]), .Y(n3412) );
  CLKINVX1 U38 ( .A(WriteData[28]), .Y(n3411) );
  CLKINVX1 U39 ( .A(WriteData[29]), .Y(n3410) );
  CLKINVX1 U40 ( .A(WriteData[30]), .Y(n3409) );
  NOR2BX1 U41 ( .AN(n80), .B(WriteReg[0]), .Y(n66) );
  NOR2BX1 U42 ( .AN(n122), .B(WriteReg[0]), .Y(n106) );
  NOR2BX1 U43 ( .AN(n100), .B(WriteReg[0]), .Y(n86) );
  NOR2X2 U44 ( .A(n3443), .B(WriteReg[1]), .Y(n53) );
  NOR2X2 U45 ( .A(n3444), .B(WriteReg[2]), .Y(n47) );
  CLKBUFX3 U46 ( .A(n3399), .Y(n3310) );
  CLKBUFX3 U47 ( .A(n3399), .Y(n3311) );
  CLKBUFX3 U48 ( .A(n3399), .Y(n3312) );
  CLKBUFX3 U49 ( .A(n3399), .Y(n3313) );
  CLKBUFX3 U50 ( .A(n3398), .Y(n3314) );
  CLKBUFX3 U51 ( .A(n3398), .Y(n3315) );
  CLKBUFX3 U52 ( .A(n3398), .Y(n3316) );
  CLKBUFX3 U53 ( .A(n3398), .Y(n3317) );
  CLKBUFX3 U54 ( .A(n3397), .Y(n3318) );
  CLKBUFX3 U55 ( .A(n3397), .Y(n3319) );
  CLKBUFX3 U56 ( .A(n3397), .Y(n3320) );
  CLKBUFX3 U57 ( .A(n3397), .Y(n3321) );
  CLKBUFX3 U58 ( .A(n3396), .Y(n3322) );
  CLKBUFX3 U59 ( .A(n3396), .Y(n3323) );
  CLKBUFX3 U60 ( .A(n3396), .Y(n3324) );
  CLKBUFX3 U61 ( .A(n3396), .Y(n3325) );
  CLKBUFX3 U62 ( .A(n3395), .Y(n3326) );
  CLKBUFX3 U63 ( .A(n3395), .Y(n3327) );
  CLKBUFX3 U64 ( .A(n3395), .Y(n3328) );
  CLKBUFX3 U65 ( .A(n3395), .Y(n3329) );
  CLKBUFX3 U66 ( .A(n3394), .Y(n3330) );
  CLKBUFX3 U67 ( .A(n3394), .Y(n3331) );
  CLKBUFX3 U68 ( .A(n3394), .Y(n3332) );
  CLKBUFX3 U69 ( .A(n3394), .Y(n3333) );
  CLKBUFX3 U70 ( .A(n3393), .Y(n3334) );
  CLKBUFX3 U71 ( .A(n3393), .Y(n3335) );
  CLKBUFX3 U72 ( .A(n3393), .Y(n3336) );
  CLKBUFX3 U73 ( .A(n3393), .Y(n3337) );
  CLKBUFX3 U74 ( .A(n3392), .Y(n3338) );
  CLKBUFX3 U75 ( .A(n3392), .Y(n3339) );
  CLKBUFX3 U76 ( .A(n3392), .Y(n3340) );
  CLKBUFX3 U77 ( .A(n3392), .Y(n3341) );
  CLKBUFX3 U78 ( .A(n3391), .Y(n3342) );
  CLKBUFX3 U79 ( .A(n3391), .Y(n3343) );
  CLKBUFX3 U80 ( .A(n3391), .Y(n3344) );
  CLKBUFX3 U81 ( .A(n3391), .Y(n3345) );
  CLKBUFX3 U82 ( .A(n3390), .Y(n3346) );
  CLKBUFX3 U83 ( .A(n3390), .Y(n3347) );
  CLKBUFX3 U84 ( .A(n3390), .Y(n3348) );
  CLKBUFX3 U85 ( .A(n3390), .Y(n3349) );
  CLKBUFX3 U86 ( .A(n3389), .Y(n3350) );
  CLKBUFX3 U87 ( .A(n3389), .Y(n3351) );
  CLKBUFX3 U88 ( .A(n3389), .Y(n3352) );
  CLKBUFX3 U89 ( .A(n3389), .Y(n3353) );
  CLKBUFX3 U90 ( .A(n3388), .Y(n3354) );
  CLKBUFX3 U91 ( .A(n3388), .Y(n3355) );
  CLKBUFX3 U92 ( .A(n3388), .Y(n3356) );
  CLKBUFX3 U93 ( .A(n3388), .Y(n3357) );
  CLKBUFX3 U94 ( .A(n3387), .Y(n3358) );
  CLKBUFX3 U95 ( .A(n3387), .Y(n3359) );
  CLKBUFX3 U96 ( .A(n3387), .Y(n3360) );
  CLKBUFX3 U97 ( .A(n3387), .Y(n3361) );
  CLKBUFX3 U98 ( .A(n3386), .Y(n3362) );
  CLKBUFX3 U99 ( .A(n3386), .Y(n3363) );
  CLKBUFX3 U100 ( .A(n3386), .Y(n3364) );
  CLKBUFX3 U101 ( .A(n3386), .Y(n3365) );
  CLKBUFX3 U102 ( .A(n3385), .Y(n3366) );
  CLKBUFX3 U103 ( .A(n3385), .Y(n3367) );
  CLKBUFX3 U104 ( .A(n3385), .Y(n3368) );
  CLKBUFX3 U105 ( .A(n3385), .Y(n3369) );
  CLKBUFX3 U106 ( .A(n3384), .Y(n3370) );
  CLKBUFX3 U107 ( .A(n3384), .Y(n3371) );
  CLKBUFX3 U108 ( .A(n3384), .Y(n3372) );
  CLKBUFX3 U109 ( .A(n3384), .Y(n3373) );
  CLKBUFX3 U110 ( .A(n3383), .Y(n3374) );
  CLKBUFX3 U111 ( .A(n3383), .Y(n3375) );
  CLKBUFX3 U112 ( .A(n3383), .Y(n3376) );
  CLKBUFX3 U113 ( .A(n3383), .Y(n3377) );
  CLKBUFX3 U114 ( .A(n3382), .Y(n3378) );
  CLKBUFX3 U115 ( .A(n3382), .Y(n3379) );
  CLKBUFX3 U116 ( .A(n3382), .Y(n3380) );
  CLKBUFX3 U117 ( .A(n3382), .Y(n3381) );
  CLKBUFX3 U118 ( .A(n3401), .Y(n3302) );
  CLKBUFX3 U119 ( .A(n3401), .Y(n3303) );
  CLKBUFX3 U120 ( .A(n3401), .Y(n3304) );
  CLKBUFX3 U121 ( .A(n3401), .Y(n3305) );
  CLKBUFX3 U122 ( .A(n3400), .Y(n3306) );
  CLKBUFX3 U123 ( .A(n3400), .Y(n3307) );
  CLKBUFX3 U124 ( .A(n3400), .Y(n3308) );
  CLKBUFX3 U125 ( .A(n3400), .Y(n3309) );
  CLKBUFX3 U126 ( .A(n3402), .Y(n3299) );
  CLKBUFX3 U127 ( .A(n3402), .Y(n3300) );
  CLKBUFX3 U128 ( .A(n3297), .Y(n3301) );
  CLKBUFX3 U129 ( .A(n3403), .Y(n3399) );
  CLKBUFX3 U130 ( .A(n3403), .Y(n3398) );
  CLKBUFX3 U131 ( .A(n3403), .Y(n3397) );
  CLKBUFX3 U132 ( .A(n3404), .Y(n3396) );
  CLKBUFX3 U133 ( .A(n3404), .Y(n3395) );
  CLKBUFX3 U134 ( .A(n3404), .Y(n3394) );
  CLKBUFX3 U135 ( .A(n3405), .Y(n3393) );
  CLKBUFX3 U136 ( .A(n3405), .Y(n3392) );
  CLKBUFX3 U137 ( .A(n3405), .Y(n3391) );
  CLKBUFX3 U138 ( .A(n3406), .Y(n3390) );
  CLKBUFX3 U139 ( .A(n3406), .Y(n3389) );
  CLKBUFX3 U140 ( .A(n3406), .Y(n3388) );
  CLKBUFX3 U141 ( .A(n3407), .Y(n3387) );
  CLKBUFX3 U142 ( .A(n3407), .Y(n3386) );
  CLKBUFX3 U143 ( .A(n3407), .Y(n3385) );
  CLKBUFX3 U144 ( .A(n3298), .Y(n3384) );
  CLKBUFX3 U145 ( .A(n3405), .Y(n3383) );
  CLKBUFX3 U146 ( .A(n3406), .Y(n3382) );
  CLKBUFX3 U147 ( .A(n3298), .Y(n3403) );
  CLKBUFX3 U148 ( .A(n3298), .Y(n3404) );
  CLKBUFX3 U149 ( .A(n3297), .Y(n3405) );
  CLKBUFX3 U150 ( .A(n3297), .Y(n3406) );
  CLKBUFX3 U151 ( .A(n3297), .Y(n3407) );
  CLKBUFX3 U152 ( .A(n3402), .Y(n3401) );
  CLKBUFX3 U153 ( .A(n3402), .Y(n3400) );
  CLKBUFX3 U154 ( .A(n3298), .Y(n3402) );
  NOR2X1 U155 ( .A(n3079), .B(n3099), .Y(n2955) );
  NOR2X1 U156 ( .A(n3079), .B(n3099), .Y(n2965) );
  NOR2X1 U157 ( .A(n3072), .B(n3099), .Y(n2970) );
  NOR2X1 U158 ( .A(n3077), .B(n3099), .Y(n2935) );
  NOR2X1 U159 ( .A(n3077), .B(n3099), .Y(n2940) );
  NOR2X1 U160 ( .A(n3077), .B(n3099), .Y(n2945) );
  NOR2X1 U161 ( .A(n3077), .B(n3099), .Y(n2950) );
  NOR2X1 U162 ( .A(n3077), .B(n3099), .Y(n2930) );
  NOR2X1 U163 ( .A(n2539), .B(n2571), .Y(n2403) );
  NOR2X1 U164 ( .A(n2549), .B(n2571), .Y(n2408) );
  NOR2X1 U165 ( .A(n2549), .B(n2571), .Y(n2413) );
  NOR2X1 U166 ( .A(n2541), .B(n2571), .Y(n2418) );
  NOR2X1 U167 ( .A(n2545), .B(n2571), .Y(n2423) );
  NOR2X1 U168 ( .A(n2539), .B(n2571), .Y(n2428) );
  NOR2X1 U169 ( .A(n2542), .B(n2571), .Y(n2438) );
  NOR2X1 U170 ( .A(n2540), .B(n2571), .Y(n2443) );
  NOR2X1 U171 ( .A(n3075), .B(n3101), .Y(n3050) );
  NOR2X1 U172 ( .A(n3075), .B(n3101), .Y(n3025) );
  NOR2X1 U173 ( .A(n2548), .B(n2573), .Y(n2498) );
  NOR2X1 U174 ( .A(n2548), .B(n2573), .Y(n2523) );
  NOR2X1 U175 ( .A(n3079), .B(n3100), .Y(n2960) );
  NOR2X1 U176 ( .A(n3077), .B(n3100), .Y(n2925) );
  NOR2X1 U177 ( .A(n3076), .B(n3101), .Y(n3035) );
  NOR2X1 U178 ( .A(n3076), .B(n3101), .Y(n3040) );
  NOR2X1 U179 ( .A(n3069), .B(n3101), .Y(n3045) );
  NOR2X1 U180 ( .A(n3076), .B(n3101), .Y(n3015) );
  NOR2X1 U181 ( .A(n3078), .B(n3101), .Y(n3020) );
  NOR2X1 U182 ( .A(n3076), .B(n3101), .Y(n3030) );
  NOR2X1 U183 ( .A(n3077), .B(n3100), .Y(n2995) );
  NOR2X1 U184 ( .A(n3076), .B(n3100), .Y(n3000) );
  NOR2X1 U185 ( .A(n3076), .B(n3100), .Y(n3005) );
  NOR2X1 U186 ( .A(n3076), .B(n3100), .Y(n3010) );
  NOR2X1 U187 ( .A(n3079), .B(n3100), .Y(n2975) );
  NOR2X1 U188 ( .A(n3079), .B(n3100), .Y(n2980) );
  NOR2X1 U189 ( .A(n3076), .B(n3100), .Y(n2985) );
  NOR2X1 U190 ( .A(n3070), .B(n3100), .Y(n2990) );
  NOR2X1 U191 ( .A(n2542), .B(n2572), .Y(n2398) );
  NOR2X1 U192 ( .A(n2541), .B(n2572), .Y(n2433) );
  NOR2X1 U193 ( .A(n2541), .B(n2572), .Y(n2448) );
  NOR2X1 U194 ( .A(n2540), .B(n2572), .Y(n2453) );
  NOR2X1 U195 ( .A(n2550), .B(n2572), .Y(n2458) );
  NOR2X1 U196 ( .A(n2550), .B(n2572), .Y(n2463) );
  NOR2X1 U197 ( .A(n2550), .B(n2572), .Y(n2468) );
  NOR2X1 U198 ( .A(n2549), .B(n2572), .Y(n2473) );
  NOR2X1 U199 ( .A(n2549), .B(n2572), .Y(n2478) );
  NOR2X1 U200 ( .A(n2549), .B(n2572), .Y(n2483) );
  NOR2X1 U201 ( .A(n2549), .B(n2573), .Y(n2488) );
  NOR2X1 U202 ( .A(n2550), .B(n2573), .Y(n2493) );
  NOR2X1 U203 ( .A(n2549), .B(n2573), .Y(n2503) );
  NOR2X1 U204 ( .A(n2549), .B(n2573), .Y(n2508) );
  NOR2X1 U205 ( .A(n2549), .B(n2573), .Y(n2513) );
  NOR2X1 U206 ( .A(n2550), .B(n2573), .Y(n2518) );
  CLKBUFX3 U207 ( .A(rst_n), .Y(n3298) );
  CLKBUFX3 U208 ( .A(rst_n), .Y(n3297) );
  CLKBUFX3 U209 ( .A(n3079), .Y(n3074) );
  CLKBUFX3 U210 ( .A(n2551), .Y(n2547) );
  CLKBUFX3 U211 ( .A(n2553), .Y(n2568) );
  CLKBUFX3 U212 ( .A(n2553), .Y(n2560) );
  CLKBUFX3 U213 ( .A(n2553), .Y(n2559) );
  CLKBUFX3 U214 ( .A(n2553), .Y(n2558) );
  CLKBUFX3 U215 ( .A(n2553), .Y(n2557) );
  CLKBUFX3 U216 ( .A(n2553), .Y(n2556) );
  CLKBUFX3 U217 ( .A(n2553), .Y(n2555) );
  CLKBUFX3 U218 ( .A(n2553), .Y(n2554) );
  CLKBUFX3 U219 ( .A(n2552), .Y(n2567) );
  CLKBUFX3 U220 ( .A(n2552), .Y(n2566) );
  CLKBUFX3 U221 ( .A(n2552), .Y(n2565) );
  CLKBUFX3 U222 ( .A(n2552), .Y(n2564) );
  CLKBUFX3 U223 ( .A(n2552), .Y(n2563) );
  CLKBUFX3 U224 ( .A(n2552), .Y(n2562) );
  CLKBUFX3 U225 ( .A(n2552), .Y(n2561) );
  CLKBUFX3 U226 ( .A(n2551), .Y(n2548) );
  CLKBUFX3 U227 ( .A(n3082), .Y(n3098) );
  CLKBUFX3 U228 ( .A(n3082), .Y(n3097) );
  CLKBUFX3 U229 ( .A(n2553), .Y(n2570) );
  CLKBUFX3 U230 ( .A(n2553), .Y(n2569) );
  CLKBUFX3 U231 ( .A(n3082), .Y(n3096) );
  NOR2X1 U232 ( .A(n2549), .B(n2573), .Y(n2373) );
  NOR2X1 U233 ( .A(n3078), .B(n3101), .Y(n2900) );
  NOR2X1 U234 ( .A(n2551), .B(n2573), .Y(n2378) );
  NOR2X1 U235 ( .A(n3078), .B(n3101), .Y(n2905) );
  NOR2X1 U236 ( .A(n2545), .B(n2573), .Y(n2383) );
  NOR2X1 U237 ( .A(n3078), .B(n3101), .Y(n2910) );
  NOR2X1 U238 ( .A(n3078), .B(n3100), .Y(n2915) );
  NOR2X1 U239 ( .A(n2548), .B(n2572), .Y(n2388) );
  CLKBUFX3 U240 ( .A(n3082), .Y(n3083) );
  CLKBUFX3 U241 ( .A(n3082), .Y(n3089) );
  CLKBUFX3 U242 ( .A(n3082), .Y(n3084) );
  CLKBUFX3 U243 ( .A(n3080), .Y(n3085) );
  CLKBUFX3 U244 ( .A(n3082), .Y(n3088) );
  CLKBUFX3 U245 ( .A(n3082), .Y(n3086) );
  CLKBUFX3 U246 ( .A(n3082), .Y(n3087) );
  CLKBUFX3 U247 ( .A(n3080), .Y(n3091) );
  CLKBUFX3 U248 ( .A(n3082), .Y(n3090) );
  CLKBUFX3 U249 ( .A(n3080), .Y(n3092) );
  CLKBUFX3 U250 ( .A(n3080), .Y(n3094) );
  CLKBUFX3 U251 ( .A(n3080), .Y(n3093) );
  CLKBUFX3 U252 ( .A(n3080), .Y(n3095) );
  BUFX4 U253 ( .A(n3079), .Y(n3065) );
  BUFX4 U254 ( .A(n2551), .Y(n2542) );
  BUFX4 U255 ( .A(n3075), .Y(n3068) );
  BUFX4 U256 ( .A(N8), .Y(n3066) );
  BUFX4 U257 ( .A(N8), .Y(n3067) );
  BUFX4 U258 ( .A(n3079), .Y(n3069) );
  BUFX4 U259 ( .A(n3079), .Y(n3070) );
  BUFX4 U260 ( .A(n3079), .Y(n3072) );
  BUFX4 U261 ( .A(n3079), .Y(n3071) );
  BUFX4 U262 ( .A(n3079), .Y(n3073) );
  BUFX4 U263 ( .A(n2551), .Y(n2541) );
  BUFX4 U264 ( .A(n2551), .Y(n2540) );
  BUFX4 U265 ( .A(n2551), .Y(n2539) );
  BUFX4 U266 ( .A(n2548), .Y(n2538) );
  BUFX4 U267 ( .A(n2551), .Y(n2546) );
  BUFX4 U268 ( .A(n2551), .Y(n2545) );
  BUFX4 U269 ( .A(n2550), .Y(n2544) );
  BUFX4 U270 ( .A(n2551), .Y(n2543) );
  CLKBUFX3 U271 ( .A(n3079), .Y(n3075) );
  CLKBUFX3 U272 ( .A(n3079), .Y(n3077) );
  CLKBUFX3 U273 ( .A(n3079), .Y(n3076) );
  CLKBUFX3 U274 ( .A(N3), .Y(n2549) );
  CLKBUFX3 U275 ( .A(n2551), .Y(n2550) );
  CLKBUFX3 U276 ( .A(n3268), .Y(n3271) );
  CLKBUFX3 U277 ( .A(n3236), .Y(n3239) );
  CLKBUFX3 U278 ( .A(n101), .Y(n3207) );
  CLKBUFX3 U279 ( .A(n3172), .Y(n3175) );
  INVX3 U280 ( .A(n3268), .Y(n3269) );
  INVX3 U281 ( .A(n3268), .Y(n3270) );
  INVX3 U282 ( .A(n3236), .Y(n3237) );
  INVX3 U283 ( .A(n3236), .Y(n3238) );
  INVX3 U284 ( .A(n101), .Y(n3205) );
  INVX3 U285 ( .A(n123), .Y(n3173) );
  INVX3 U286 ( .A(n3172), .Y(n3174) );
  INVX3 U287 ( .A(n101), .Y(n3206) );
  CLKBUFX3 U288 ( .A(N2), .Y(n2553) );
  CLKBUFX3 U289 ( .A(n3056), .Y(n3060) );
  CLKBUFX3 U290 ( .A(n3056), .Y(n3059) );
  CLKBUFX3 U291 ( .A(n3056), .Y(n3057) );
  CLKBUFX3 U292 ( .A(n3056), .Y(n3058) );
  CLKBUFX3 U293 ( .A(N5), .Y(n2533) );
  CLKBUFX3 U294 ( .A(n2529), .Y(n2532) );
  CLKBUFX3 U295 ( .A(n2529), .Y(n2531) );
  CLKBUFX3 U296 ( .A(n2529), .Y(n2530) );
  CLKBUFX3 U297 ( .A(n3079), .Y(n3078) );
  CLKBUFX3 U298 ( .A(n3061), .Y(n3064) );
  CLKBUFX3 U299 ( .A(n3061), .Y(n3062) );
  CLKBUFX3 U300 ( .A(n3061), .Y(n3063) );
  CLKBUFX3 U301 ( .A(n2534), .Y(n2537) );
  CLKBUFX3 U302 ( .A(n2534), .Y(n2536) );
  CLKBUFX3 U303 ( .A(n2534), .Y(n2535) );
  CLKBUFX3 U304 ( .A(n3080), .Y(n3081) );
  CLKBUFX3 U305 ( .A(N7), .Y(n3082) );
  CLKBUFX3 U306 ( .A(N9), .Y(n3061) );
  CLKBUFX3 U307 ( .A(n3296), .Y(n3294) );
  CLKBUFX3 U308 ( .A(n3296), .Y(n3295) );
  CLKBUFX3 U309 ( .A(n3288), .Y(n3291) );
  CLKBUFX3 U310 ( .A(n3284), .Y(n3287) );
  CLKBUFX3 U311 ( .A(n51), .Y(n3283) );
  CLKBUFX3 U312 ( .A(n3276), .Y(n3279) );
  CLKBUFX3 U313 ( .A(n56), .Y(n3275) );
  CLKBUFX3 U314 ( .A(n3264), .Y(n3267) );
  CLKBUFX3 U315 ( .A(n3260), .Y(n3263) );
  CLKBUFX3 U316 ( .A(n3256), .Y(n3259) );
  CLKBUFX3 U317 ( .A(n3252), .Y(n3255) );
  CLKBUFX3 U318 ( .A(n3248), .Y(n3251) );
  CLKBUFX3 U319 ( .A(n3244), .Y(n3247) );
  CLKBUFX3 U320 ( .A(n3240), .Y(n3243) );
  CLKBUFX3 U321 ( .A(n84), .Y(n3235) );
  CLKBUFX3 U322 ( .A(n87), .Y(n3231) );
  CLKBUFX3 U323 ( .A(n90), .Y(n3227) );
  CLKBUFX3 U324 ( .A(n92), .Y(n3223) );
  CLKBUFX3 U325 ( .A(n3216), .Y(n3219) );
  CLKBUFX3 U326 ( .A(n3200), .Y(n3203) );
  CLKBUFX3 U327 ( .A(n3196), .Y(n3199) );
  CLKBUFX3 U328 ( .A(n3192), .Y(n3195) );
  CLKBUFX3 U329 ( .A(n3188), .Y(n3191) );
  CLKBUFX3 U330 ( .A(n3184), .Y(n3187) );
  CLKBUFX3 U331 ( .A(n3180), .Y(n3183) );
  CLKBUFX3 U332 ( .A(n3176), .Y(n3179) );
  INVX3 U333 ( .A(n45), .Y(n3289) );
  INVX3 U334 ( .A(n3284), .Y(n3285) );
  INVX3 U335 ( .A(n51), .Y(n3281) );
  INVX3 U336 ( .A(n3280), .Y(n3282) );
  INVX3 U337 ( .A(n3276), .Y(n3277) );
  INVX3 U338 ( .A(n3276), .Y(n3278) );
  INVX3 U339 ( .A(n56), .Y(n3273) );
  INVX3 U340 ( .A(n3272), .Y(n3274) );
  INVX3 U341 ( .A(n3264), .Y(n3265) );
  INVX3 U342 ( .A(n3264), .Y(n3266) );
  INVX3 U343 ( .A(n3260), .Y(n3261) );
  INVX3 U344 ( .A(n3260), .Y(n3262) );
  INVX3 U345 ( .A(n3256), .Y(n3257) );
  INVX3 U346 ( .A(n3256), .Y(n3258) );
  INVX3 U347 ( .A(n3252), .Y(n3253) );
  INVX3 U348 ( .A(n3252), .Y(n3254) );
  INVX3 U349 ( .A(n3248), .Y(n3249) );
  INVX3 U350 ( .A(n3248), .Y(n3250) );
  INVX3 U351 ( .A(n3244), .Y(n3245) );
  INVX3 U352 ( .A(n3244), .Y(n3246) );
  INVX3 U353 ( .A(n3240), .Y(n3241) );
  INVX3 U354 ( .A(n3240), .Y(n3242) );
  INVX3 U355 ( .A(n84), .Y(n3233) );
  INVX3 U356 ( .A(n3232), .Y(n3234) );
  INVX3 U357 ( .A(n87), .Y(n3229) );
  INVX3 U358 ( .A(n3228), .Y(n3230) );
  INVX3 U359 ( .A(n90), .Y(n3225) );
  INVX3 U360 ( .A(n3224), .Y(n3226) );
  INVX3 U361 ( .A(n92), .Y(n3221) );
  INVX3 U362 ( .A(n3220), .Y(n3222) );
  INVX3 U363 ( .A(n3216), .Y(n3217) );
  INVX3 U364 ( .A(n96), .Y(n3214) );
  INVX3 U365 ( .A(n96), .Y(n3215) );
  INVX3 U366 ( .A(n98), .Y(n3210) );
  INVX3 U367 ( .A(n98), .Y(n3211) );
  INVX3 U368 ( .A(n3200), .Y(n3201) );
  INVX3 U369 ( .A(n3200), .Y(n3202) );
  INVX3 U370 ( .A(n107), .Y(n3197) );
  INVX3 U371 ( .A(n3196), .Y(n3198) );
  INVX3 U372 ( .A(n3192), .Y(n3193) );
  INVX3 U373 ( .A(n3192), .Y(n3194) );
  INVX3 U374 ( .A(n112), .Y(n3189) );
  INVX3 U375 ( .A(n3188), .Y(n3190) );
  INVX3 U376 ( .A(n3184), .Y(n3185) );
  INVX3 U377 ( .A(n3184), .Y(n3186) );
  INVX3 U378 ( .A(n117), .Y(n3181) );
  INVX3 U379 ( .A(n3180), .Y(n3182) );
  INVX3 U380 ( .A(n3176), .Y(n3177) );
  INVX3 U381 ( .A(n3176), .Y(n3178) );
  INVX3 U382 ( .A(n3296), .Y(n3293) );
  INVX3 U383 ( .A(n3288), .Y(n3290) );
  INVX3 U384 ( .A(n3284), .Y(n3286) );
  INVX3 U385 ( .A(n3216), .Y(n3218) );
  CLKBUFX3 U386 ( .A(n60), .Y(n3268) );
  CLKBUFX3 U387 ( .A(n81), .Y(n3236) );
  CLKBUFX3 U388 ( .A(n101), .Y(n3204) );
  CLKBUFX3 U389 ( .A(n123), .Y(n3172) );
  CLKBUFX3 U390 ( .A(n3439), .Y(n3164) );
  CLKBUFX3 U391 ( .A(n3438), .Y(n3162) );
  CLKBUFX3 U392 ( .A(n3437), .Y(n3160) );
  CLKBUFX3 U393 ( .A(n3436), .Y(n3158) );
  CLKBUFX3 U394 ( .A(n3435), .Y(n3156) );
  CLKBUFX3 U395 ( .A(n3434), .Y(n3154) );
  CLKBUFX3 U396 ( .A(n3433), .Y(n3152) );
  CLKBUFX3 U397 ( .A(n3432), .Y(n3150) );
  CLKBUFX3 U398 ( .A(n3431), .Y(n3148) );
  CLKBUFX3 U399 ( .A(n3430), .Y(n3146) );
  CLKBUFX3 U400 ( .A(n3429), .Y(n3144) );
  CLKBUFX3 U401 ( .A(n3428), .Y(n3142) );
  CLKBUFX3 U402 ( .A(n3427), .Y(n3140) );
  CLKBUFX3 U403 ( .A(n3426), .Y(n3138) );
  CLKBUFX3 U404 ( .A(n3425), .Y(n3136) );
  CLKBUFX3 U405 ( .A(n3424), .Y(n3134) );
  CLKBUFX3 U406 ( .A(n3423), .Y(n3132) );
  CLKBUFX3 U407 ( .A(n3422), .Y(n3130) );
  CLKBUFX3 U408 ( .A(n3421), .Y(n3128) );
  CLKBUFX3 U409 ( .A(n3420), .Y(n3126) );
  CLKBUFX3 U410 ( .A(n3419), .Y(n3124) );
  CLKBUFX3 U411 ( .A(n3418), .Y(n3122) );
  CLKBUFX3 U412 ( .A(n3417), .Y(n3120) );
  CLKBUFX3 U413 ( .A(n3416), .Y(n3118) );
  CLKBUFX3 U414 ( .A(n3415), .Y(n3116) );
  CLKBUFX3 U415 ( .A(n3414), .Y(n3114) );
  CLKBUFX3 U416 ( .A(n3413), .Y(n3112) );
  CLKBUFX3 U417 ( .A(n3412), .Y(n3110) );
  CLKBUFX3 U418 ( .A(n3411), .Y(n3108) );
  CLKBUFX3 U419 ( .A(n3410), .Y(n3106) );
  CLKBUFX3 U420 ( .A(n3409), .Y(n3104) );
  CLKBUFX3 U421 ( .A(n3408), .Y(n3102) );
  CLKBUFX3 U422 ( .A(N11), .Y(n3055) );
  CLKBUFX3 U423 ( .A(N11), .Y(n3054) );
  CLKBUFX3 U424 ( .A(n2528), .Y(n2527) );
  CLKBUFX3 U425 ( .A(n125), .Y(n3170) );
  CLKBUFX3 U426 ( .A(n132), .Y(n3167) );
  CLKBUFX3 U427 ( .A(n125), .Y(n3171) );
  CLKBUFX3 U428 ( .A(n132), .Y(n3168) );
  CLKBUFX3 U429 ( .A(n125), .Y(n3169) );
  CLKBUFX3 U430 ( .A(n132), .Y(n3166) );
  CLKBUFX3 U431 ( .A(N7), .Y(n3080) );
  CLKBUFX3 U432 ( .A(N2), .Y(n2552) );
  CLKBUFX3 U433 ( .A(N10), .Y(n3056) );
  CLKBUFX3 U434 ( .A(N4), .Y(n2534) );
  CLKBUFX3 U435 ( .A(N5), .Y(n2529) );
  CLKBUFX3 U436 ( .A(n3439), .Y(n3165) );
  CLKBUFX3 U437 ( .A(n3438), .Y(n3163) );
  CLKBUFX3 U438 ( .A(n3437), .Y(n3161) );
  CLKBUFX3 U439 ( .A(n3436), .Y(n3159) );
  CLKBUFX3 U440 ( .A(n3435), .Y(n3157) );
  CLKBUFX3 U441 ( .A(n3434), .Y(n3155) );
  CLKBUFX3 U442 ( .A(n3433), .Y(n3153) );
  CLKBUFX3 U443 ( .A(n3432), .Y(n3151) );
  CLKBUFX3 U444 ( .A(n3431), .Y(n3149) );
  CLKBUFX3 U445 ( .A(n3430), .Y(n3147) );
  CLKBUFX3 U446 ( .A(n3429), .Y(n3145) );
  CLKBUFX3 U447 ( .A(n3428), .Y(n3143) );
  CLKBUFX3 U448 ( .A(n3427), .Y(n3141) );
  CLKBUFX3 U449 ( .A(n3426), .Y(n3139) );
  CLKBUFX3 U450 ( .A(n3425), .Y(n3137) );
  CLKBUFX3 U451 ( .A(n3424), .Y(n3135) );
  CLKBUFX3 U452 ( .A(n3423), .Y(n3133) );
  CLKBUFX3 U453 ( .A(n3422), .Y(n3131) );
  CLKBUFX3 U454 ( .A(n3421), .Y(n3129) );
  CLKBUFX3 U455 ( .A(n3420), .Y(n3127) );
  CLKBUFX3 U456 ( .A(n3419), .Y(n3125) );
  CLKBUFX3 U457 ( .A(n3418), .Y(n3123) );
  CLKBUFX3 U458 ( .A(n3417), .Y(n3121) );
  CLKBUFX3 U459 ( .A(n3416), .Y(n3119) );
  CLKBUFX3 U460 ( .A(n3415), .Y(n3117) );
  CLKBUFX3 U461 ( .A(n3414), .Y(n3115) );
  CLKBUFX3 U462 ( .A(n3413), .Y(n3113) );
  CLKBUFX3 U463 ( .A(n3412), .Y(n3111) );
  CLKBUFX3 U464 ( .A(n3411), .Y(n3109) );
  CLKBUFX3 U465 ( .A(n3410), .Y(n3107) );
  CLKBUFX3 U466 ( .A(n3409), .Y(n3105) );
  CLKBUFX3 U467 ( .A(n3408), .Y(n3103) );
  CLKBUFX3 U468 ( .A(n45), .Y(n3288) );
  CLKBUFX3 U469 ( .A(n49), .Y(n3284) );
  CLKBUFX3 U470 ( .A(n51), .Y(n3280) );
  CLKBUFX3 U471 ( .A(n54), .Y(n3276) );
  CLKBUFX3 U472 ( .A(n56), .Y(n3272) );
  CLKBUFX3 U473 ( .A(n64), .Y(n3264) );
  CLKBUFX3 U474 ( .A(n67), .Y(n3260) );
  CLKBUFX3 U475 ( .A(n70), .Y(n3256) );
  CLKBUFX3 U476 ( .A(n72), .Y(n3252) );
  CLKBUFX3 U477 ( .A(n74), .Y(n3248) );
  CLKBUFX3 U478 ( .A(n76), .Y(n3244) );
  CLKBUFX3 U479 ( .A(n78), .Y(n3240) );
  CLKBUFX3 U480 ( .A(n84), .Y(n3232) );
  CLKBUFX3 U481 ( .A(n87), .Y(n3228) );
  CLKBUFX3 U482 ( .A(n90), .Y(n3224) );
  CLKBUFX3 U483 ( .A(n92), .Y(n3220) );
  CLKBUFX3 U484 ( .A(n96), .Y(n3212) );
  CLKBUFX3 U485 ( .A(n96), .Y(n3213) );
  CLKBUFX3 U486 ( .A(n98), .Y(n3208) );
  CLKBUFX3 U487 ( .A(n98), .Y(n3209) );
  CLKBUFX3 U488 ( .A(n104), .Y(n3200) );
  CLKBUFX3 U489 ( .A(n107), .Y(n3196) );
  CLKBUFX3 U490 ( .A(n110), .Y(n3192) );
  CLKBUFX3 U491 ( .A(n112), .Y(n3188) );
  CLKBUFX3 U492 ( .A(n115), .Y(n3184) );
  CLKBUFX3 U493 ( .A(n117), .Y(n3180) );
  CLKBUFX3 U494 ( .A(n120), .Y(n3176) );
  CLKINVX1 U495 ( .A(n3292), .Y(n3296) );
  NAND2X1 U496 ( .A(n58), .B(n44), .Y(n60) );
  NAND2X1 U497 ( .A(n69), .B(n58), .Y(n81) );
  NAND2X1 U498 ( .A(n89), .B(n58), .Y(n101) );
  NAND2X1 U499 ( .A(n109), .B(n58), .Y(n123) );
  OAI2BB2XL U500 ( .B0(n3104), .B1(n3167), .A0N(prev_ReadData1[30]), .A1N(
        n3167), .Y(ReadData1[30]) );
  MXI2X1 U501 ( .A(n91), .B(n93), .S0(n2527), .Y(prev_ReadData1[30]) );
  MX4X1 U502 ( .A(n2354), .B(n2352), .C(n2353), .D(n2351), .S0(n2533), .S1(
        n2537), .Y(n93) );
  OAI2BB2XL U503 ( .B0(n3146), .B1(n3167), .A0N(prev_ReadData1[9]), .A1N(n3166), .Y(ReadData1[9]) );
  MXI2X1 U504 ( .A(n20), .B(n21), .S0(n2528), .Y(prev_ReadData1[9]) );
  MX4X1 U505 ( .A(n2190), .B(n2188), .C(n2189), .D(n2187), .S0(n2530), .S1(
        n2534), .Y(n20) );
  OAI2BB2XL U506 ( .B0(n3150), .B1(n3167), .A0N(prev_ReadData1[7]), .A1N(n3168), .Y(ReadData1[7]) );
  MXI2X1 U507 ( .A(n16), .B(n17), .S0(n2528), .Y(prev_ReadData1[7]) );
  MX4X1 U508 ( .A(n2174), .B(n2172), .C(n2173), .D(n2171), .S0(n2529), .S1(
        n2534), .Y(n16) );
  OAI2BB2XL U509 ( .B0(n3152), .B1(n3167), .A0N(prev_ReadData1[6]), .A1N(n3168), .Y(ReadData1[6]) );
  MXI2X1 U510 ( .A(n14), .B(n15), .S0(n2528), .Y(prev_ReadData1[6]) );
  MX4X1 U511 ( .A(n2166), .B(n2164), .C(n2165), .D(n2163), .S0(n2529), .S1(
        n2536), .Y(n14) );
  OAI2BB2XL U512 ( .B0(n3154), .B1(n3167), .A0N(prev_ReadData1[5]), .A1N(n3168), .Y(ReadData1[5]) );
  MXI2X1 U513 ( .A(n12), .B(n13), .S0(n2528), .Y(prev_ReadData1[5]) );
  MX4X1 U514 ( .A(n2158), .B(n2156), .C(n2157), .D(n2155), .S0(n2529), .S1(
        n2537), .Y(n12) );
  OAI2BB2XL U515 ( .B0(n3158), .B1(n3167), .A0N(prev_ReadData1[3]), .A1N(n3168), .Y(ReadData1[3]) );
  MXI2X1 U516 ( .A(n7), .B(n8), .S0(n2528), .Y(prev_ReadData1[3]) );
  MX4X1 U517 ( .A(n2142), .B(n2140), .C(n2141), .D(n2139), .S0(n2529), .S1(
        n2537), .Y(n7) );
  OAI2BB2XL U518 ( .B0(n3126), .B1(n3169), .A0N(prev_ReadData2[19]), .A1N(
        n3171), .Y(ReadData2[19]) );
  MXI2X1 U519 ( .A(n2612), .B(n2613), .S0(n3054), .Y(prev_ReadData2[19]) );
  MX4X1 U520 ( .A(n2793), .B(n2791), .C(n2792), .D(n2790), .S0(N10), .S1(n3063), .Y(n2613) );
  OAI2BB2XL U521 ( .B0(n3102), .B1(n3167), .A0N(prev_ReadData1[31]), .A1N(
        n3168), .Y(ReadData1[31]) );
  MXI2X1 U522 ( .A(n95), .B(n97), .S0(n2527), .Y(prev_ReadData1[31]) );
  MX4X1 U523 ( .A(n2362), .B(n2360), .C(n2361), .D(n2359), .S0(n2533), .S1(
        n2537), .Y(n97) );
  OAI2BB2XL U524 ( .B0(n3106), .B1(n132), .A0N(prev_ReadData1[29]), .A1N(n3167), .Y(ReadData1[29]) );
  MXI2X1 U525 ( .A(n85), .B(n88), .S0(n2527), .Y(prev_ReadData1[29]) );
  MX4X1 U526 ( .A(n2346), .B(n2344), .C(n2345), .D(n2343), .S0(n2533), .S1(
        n2537), .Y(n88) );
  OAI2BB2XL U527 ( .B0(n3110), .B1(n3166), .A0N(prev_ReadData1[27]), .A1N(
        n3167), .Y(ReadData1[27]) );
  MXI2X1 U528 ( .A(n77), .B(n79), .S0(n2527), .Y(prev_ReadData1[27]) );
  MX4X1 U529 ( .A(n2330), .B(n2328), .C(n2329), .D(n2327), .S0(n2533), .S1(
        n2537), .Y(n79) );
  OAI2BB2XL U530 ( .B0(n3112), .B1(n3166), .A0N(prev_ReadData1[26]), .A1N(
        n3167), .Y(ReadData1[26]) );
  MXI2X1 U531 ( .A(n73), .B(n75), .S0(n2527), .Y(prev_ReadData1[26]) );
  MX4X1 U532 ( .A(n2322), .B(n2320), .C(n2321), .D(n2319), .S0(n2533), .S1(
        n2537), .Y(n75) );
  OAI2BB2XL U533 ( .B0(n3114), .B1(n132), .A0N(prev_ReadData1[25]), .A1N(n3167), .Y(ReadData1[25]) );
  MXI2X1 U534 ( .A(n68), .B(n71), .S0(n2527), .Y(prev_ReadData1[25]) );
  MX4X1 U535 ( .A(n2314), .B(n2312), .C(n2313), .D(n2311), .S0(n2532), .S1(
        n2536), .Y(n71) );
  OAI2BB2XL U536 ( .B0(n3118), .B1(n3167), .A0N(prev_ReadData1[23]), .A1N(
        n3167), .Y(ReadData1[23]) );
  MXI2X1 U537 ( .A(n61), .B(n62), .S0(n2527), .Y(prev_ReadData1[23]) );
  MX4X1 U538 ( .A(n2298), .B(n2296), .C(n2297), .D(n2295), .S0(n2532), .S1(
        n2536), .Y(n62) );
  OAI2BB2XL U539 ( .B0(n3120), .B1(n132), .A0N(prev_ReadData1[22]), .A1N(n3168), .Y(ReadData1[22]) );
  MXI2X1 U540 ( .A(n55), .B(n57), .S0(n2527), .Y(prev_ReadData1[22]) );
  MX4X1 U541 ( .A(n2290), .B(n2288), .C(n2289), .D(n2287), .S0(n2532), .S1(
        n2536), .Y(n57) );
  OAI2BB2XL U542 ( .B0(n3122), .B1(n3167), .A0N(prev_ReadData1[21]), .A1N(
        n3168), .Y(ReadData1[21]) );
  MXI2X1 U543 ( .A(n50), .B(n52), .S0(n2527), .Y(prev_ReadData1[21]) );
  MX4X1 U544 ( .A(n2282), .B(n2280), .C(n2281), .D(n2279), .S0(n2532), .S1(
        n2536), .Y(n52) );
  OAI2BB2XL U545 ( .B0(n3126), .B1(n3166), .A0N(prev_ReadData1[19]), .A1N(
        n3168), .Y(ReadData1[19]) );
  MXI2X1 U546 ( .A(n40), .B(n41), .S0(n2528), .Y(prev_ReadData1[19]) );
  MX4X1 U547 ( .A(n2266), .B(n2264), .C(n2265), .D(n2263), .S0(n2531), .S1(
        n2535), .Y(n41) );
  OAI2BB2XL U548 ( .B0(n3128), .B1(n3166), .A0N(prev_ReadData1[18]), .A1N(
        n3168), .Y(ReadData1[18]) );
  MXI2X1 U549 ( .A(n38), .B(n39), .S0(n2528), .Y(prev_ReadData1[18]) );
  MX4X1 U550 ( .A(n2258), .B(n2256), .C(n2257), .D(n2255), .S0(n2531), .S1(
        n2535), .Y(n39) );
  OAI2BB2XL U551 ( .B0(n3130), .B1(n3166), .A0N(prev_ReadData1[17]), .A1N(
        n3168), .Y(ReadData1[17]) );
  MXI2X1 U552 ( .A(n36), .B(n37), .S0(n2528), .Y(prev_ReadData1[17]) );
  MX4X1 U553 ( .A(n2250), .B(n2248), .C(n2249), .D(n2247), .S0(n2531), .S1(
        n2535), .Y(n37) );
  OAI2BB2XL U554 ( .B0(n3134), .B1(n3166), .A0N(prev_ReadData1[15]), .A1N(
        n3168), .Y(ReadData1[15]) );
  MXI2X1 U555 ( .A(n32), .B(n33), .S0(n2528), .Y(prev_ReadData1[15]) );
  MX4X1 U556 ( .A(n2238), .B(n2236), .C(n2237), .D(n2235), .S0(n2531), .S1(
        n2535), .Y(n32) );
  OAI2BB2XL U557 ( .B0(n3136), .B1(n3166), .A0N(prev_ReadData1[14]), .A1N(
        n3168), .Y(ReadData1[14]) );
  MXI2X1 U558 ( .A(n30), .B(n31), .S0(n2528), .Y(prev_ReadData1[14]) );
  MX4X1 U559 ( .A(n2230), .B(n2228), .C(n2229), .D(n2227), .S0(n2531), .S1(
        n2535), .Y(n30) );
  OAI2BB2XL U560 ( .B0(n3138), .B1(n3166), .A0N(prev_ReadData1[13]), .A1N(
        n3166), .Y(ReadData1[13]) );
  MXI2X1 U561 ( .A(n28), .B(n29), .S0(n2528), .Y(prev_ReadData1[13]) );
  MX4X1 U562 ( .A(n2222), .B(n2220), .C(n2221), .D(n2219), .S0(n2530), .S1(
        n2534), .Y(n28) );
  OAI2BB2XL U563 ( .B0(n3142), .B1(n3166), .A0N(prev_ReadData1[11]), .A1N(
        n3168), .Y(ReadData1[11]) );
  MXI2X1 U564 ( .A(n24), .B(n25), .S0(n2528), .Y(prev_ReadData1[11]) );
  MX4X1 U565 ( .A(n2206), .B(n2204), .C(n2205), .D(n2203), .S0(n2530), .S1(
        n2537), .Y(n24) );
  OAI2BB2XL U566 ( .B0(n3144), .B1(n3166), .A0N(prev_ReadData1[10]), .A1N(
        n3168), .Y(ReadData1[10]) );
  MXI2X1 U567 ( .A(n22), .B(n23), .S0(n2528), .Y(prev_ReadData1[10]) );
  MX4X1 U568 ( .A(n2198), .B(n2196), .C(n2197), .D(n2195), .S0(n2530), .S1(
        n2534), .Y(n22) );
  OAI2BB2XL U569 ( .B0(n3160), .B1(n132), .A0N(prev_ReadData1[2]), .A1N(n3168), 
        .Y(ReadData1[2]) );
  MXI2X1 U570 ( .A(n5), .B(n6), .S0(n2528), .Y(prev_ReadData1[2]) );
  MX4X1 U571 ( .A(n2134), .B(n2132), .C(n2133), .D(n2131), .S0(n2529), .S1(
        n2535), .Y(n5) );
  OAI2BB2XL U572 ( .B0(n3162), .B1(n3166), .A0N(prev_ReadData1[1]), .A1N(n3168), .Y(ReadData1[1]) );
  MXI2X1 U573 ( .A(n3), .B(n4), .S0(n2528), .Y(prev_ReadData1[1]) );
  MX4X1 U574 ( .A(n2126), .B(n2124), .C(n2125), .D(n2123), .S0(n2532), .S1(
        n2536), .Y(n3) );
  OAI2BB2XL U575 ( .B0(n3164), .B1(n3166), .A0N(prev_ReadData1[0]), .A1N(n3168), .Y(ReadData1[0]) );
  MXI2X1 U576 ( .A(n1), .B(n2), .S0(n2527), .Y(prev_ReadData1[0]) );
  MX4X1 U577 ( .A(n108), .B(n102), .C(n105), .D(n99), .S0(n2531), .S1(n2534), 
        .Y(n2) );
  CLKBUFX3 U578 ( .A(N8), .Y(n3079) );
  CLKBUFX3 U579 ( .A(N3), .Y(n2551) );
  OAI2BB2XL U580 ( .B0(n3104), .B1(n3170), .A0N(prev_ReadData2[30]), .A1N(
        n3170), .Y(ReadData2[30]) );
  MXI2X1 U581 ( .A(n2634), .B(n2635), .S0(n3055), .Y(prev_ReadData2[30]) );
  MX4X1 U582 ( .A(n2881), .B(n2879), .C(n2880), .D(n2878), .S0(n3060), .S1(
        n3063), .Y(n2635) );
  OAI2BB2XL U583 ( .B0(n3158), .B1(n3170), .A0N(prev_ReadData2[3]), .A1N(n3171), .Y(ReadData2[3]) );
  MXI2X1 U584 ( .A(n2580), .B(n2581), .S0(n3055), .Y(prev_ReadData2[3]) );
  MX4X1 U585 ( .A(n2669), .B(n2667), .C(n2668), .D(n2666), .S0(n3057), .S1(
        n3062), .Y(n2580) );
  OAI2BB2XL U586 ( .B0(n3150), .B1(n3170), .A0N(prev_ReadData2[7]), .A1N(n3171), .Y(ReadData2[7]) );
  MXI2X1 U587 ( .A(n2588), .B(n2589), .S0(n3054), .Y(prev_ReadData2[7]) );
  MX4X1 U588 ( .A(n2701), .B(n2699), .C(n2700), .D(n2698), .S0(n3057), .S1(
        n3062), .Y(n2588) );
  OAI2BB2XL U589 ( .B0(n3152), .B1(n3170), .A0N(prev_ReadData2[6]), .A1N(n3171), .Y(ReadData2[6]) );
  MXI2X1 U590 ( .A(n2586), .B(n2587), .S0(n3054), .Y(prev_ReadData2[6]) );
  MX4X1 U591 ( .A(n2693), .B(n2691), .C(n2692), .D(n2690), .S0(n3057), .S1(
        n3062), .Y(n2586) );
  OAI2BB2XL U592 ( .B0(n3154), .B1(n3170), .A0N(prev_ReadData2[5]), .A1N(n3171), .Y(ReadData2[5]) );
  MXI2X1 U593 ( .A(n2584), .B(n2585), .S0(n3054), .Y(prev_ReadData2[5]) );
  MX4X1 U594 ( .A(n2685), .B(n2683), .C(n2684), .D(n2682), .S0(n3057), .S1(
        n3062), .Y(n2584) );
  OAI2BB2XL U595 ( .B0(n3156), .B1(n3170), .A0N(prev_ReadData2[4]), .A1N(n3171), .Y(ReadData2[4]) );
  MXI2X1 U596 ( .A(n2582), .B(n2583), .S0(n3054), .Y(prev_ReadData2[4]) );
  MX4X1 U597 ( .A(n2677), .B(n2675), .C(n2676), .D(n2674), .S0(n3057), .S1(
        n3062), .Y(n2582) );
  OAI2BB2XL U598 ( .B0(n3146), .B1(n3170), .A0N(prev_ReadData2[9]), .A1N(n3169), .Y(ReadData2[9]) );
  MXI2X1 U599 ( .A(n2592), .B(n2593), .S0(n3054), .Y(prev_ReadData2[9]) );
  MX4X1 U600 ( .A(n2717), .B(n2715), .C(n2716), .D(n2714), .S0(n3058), .S1(
        n3061), .Y(n2592) );
  OAI2BB2XL U601 ( .B0(n3148), .B1(n3170), .A0N(prev_ReadData2[8]), .A1N(n3169), .Y(ReadData2[8]) );
  MXI2X1 U602 ( .A(n2590), .B(n2591), .S0(n3054), .Y(prev_ReadData2[8]) );
  MX4X1 U603 ( .A(n2709), .B(n2707), .C(n2708), .D(n2706), .S0(n3058), .S1(
        n3063), .Y(n2590) );
  OAI2BB2XL U604 ( .B0(n3148), .B1(n3167), .A0N(prev_ReadData1[8]), .A1N(n3166), .Y(ReadData1[8]) );
  MXI2X1 U605 ( .A(n18), .B(n19), .S0(N6), .Y(prev_ReadData1[8]) );
  MX4X1 U606 ( .A(n2182), .B(n2180), .C(n2181), .D(n2179), .S0(n2530), .S1(
        n2534), .Y(n18) );
  OAI2BB2XL U607 ( .B0(n3156), .B1(n3167), .A0N(prev_ReadData1[4]), .A1N(n3168), .Y(ReadData1[4]) );
  MXI2X1 U608 ( .A(n10), .B(n11), .S0(n2528), .Y(prev_ReadData1[4]) );
  MX4X1 U609 ( .A(n2150), .B(n2148), .C(n2149), .D(n2147), .S0(N5), .S1(n2536), 
        .Y(n10) );
  OAI2BB2XL U610 ( .B0(n3128), .B1(n3169), .A0N(prev_ReadData2[18]), .A1N(
        n3171), .Y(ReadData2[18]) );
  MXI2X1 U611 ( .A(n2610), .B(n2611), .S0(n3054), .Y(prev_ReadData2[18]) );
  MX4X1 U612 ( .A(n2785), .B(n2783), .C(n2784), .D(n2782), .S0(n3056), .S1(
        n3063), .Y(n2611) );
  OAI2BB2XL U613 ( .B0(n3130), .B1(n3169), .A0N(prev_ReadData2[17]), .A1N(
        n3171), .Y(ReadData2[17]) );
  MXI2X1 U614 ( .A(n2608), .B(n2609), .S0(n3054), .Y(prev_ReadData2[17]) );
  MX4X1 U615 ( .A(n2777), .B(n2775), .C(n2776), .D(n2774), .S0(n3056), .S1(
        n3063), .Y(n2609) );
  OAI2BB2XL U616 ( .B0(n3132), .B1(n3169), .A0N(prev_ReadData2[16]), .A1N(
        n3171), .Y(ReadData2[16]) );
  MXI2X1 U617 ( .A(n2606), .B(n2607), .S0(n3054), .Y(prev_ReadData2[16]) );
  MX4X1 U618 ( .A(n2769), .B(n2767), .C(n2768), .D(n2766), .S0(n3056), .S1(
        n3063), .Y(n2607) );
  OAI2BB2XL U619 ( .B0(n3102), .B1(n3170), .A0N(prev_ReadData2[31]), .A1N(
        n3171), .Y(ReadData2[31]) );
  MXI2X1 U620 ( .A(n2636), .B(n2637), .S0(n3055), .Y(prev_ReadData2[31]) );
  MX4X1 U621 ( .A(n2889), .B(n2887), .C(n2888), .D(n2886), .S0(n3060), .S1(
        n3064), .Y(n2637) );
  OAI2BB2XL U622 ( .B0(n3106), .B1(n125), .A0N(prev_ReadData2[29]), .A1N(n3170), .Y(ReadData2[29]) );
  MXI2X1 U623 ( .A(n2632), .B(n2633), .S0(n3055), .Y(prev_ReadData2[29]) );
  MX4X1 U624 ( .A(n2873), .B(n2871), .C(n2872), .D(n2870), .S0(n3060), .S1(
        n3062), .Y(n2633) );
  OAI2BB2XL U625 ( .B0(n3108), .B1(n3166), .A0N(prev_ReadData1[28]), .A1N(
        n3167), .Y(ReadData1[28]) );
  MXI2X1 U626 ( .A(n82), .B(n83), .S0(n2527), .Y(prev_ReadData1[28]) );
  MX4X1 U627 ( .A(n2338), .B(n2336), .C(n2337), .D(n2335), .S0(n2533), .S1(
        n2537), .Y(n83) );
  OAI2BB2XL U628 ( .B0(n3108), .B1(n3169), .A0N(prev_ReadData2[28]), .A1N(
        n3170), .Y(ReadData2[28]) );
  MXI2X1 U629 ( .A(n2630), .B(n2631), .S0(n3055), .Y(prev_ReadData2[28]) );
  MX4X1 U630 ( .A(n2865), .B(n2863), .C(n2864), .D(n2862), .S0(n3060), .S1(
        n3062), .Y(n2631) );
  OAI2BB2XL U631 ( .B0(n3118), .B1(n3170), .A0N(prev_ReadData2[23]), .A1N(
        n3170), .Y(ReadData2[23]) );
  MXI2X1 U632 ( .A(n2620), .B(n2621), .S0(n3055), .Y(prev_ReadData2[23]) );
  MX4X1 U633 ( .A(n2825), .B(n2823), .C(n2824), .D(n2822), .S0(n3059), .S1(
        n3064), .Y(n2621) );
  OAI2BB2XL U634 ( .B0(n3120), .B1(n125), .A0N(prev_ReadData2[22]), .A1N(n3171), .Y(ReadData2[22]) );
  MXI2X1 U635 ( .A(n2618), .B(n2619), .S0(n3055), .Y(prev_ReadData2[22]) );
  MX4X1 U636 ( .A(n2817), .B(n2815), .C(n2816), .D(n2814), .S0(n3059), .S1(
        n3064), .Y(n2619) );
  OAI2BB2XL U637 ( .B0(n3122), .B1(n3170), .A0N(prev_ReadData2[21]), .A1N(
        n3171), .Y(ReadData2[21]) );
  MXI2X1 U638 ( .A(n2616), .B(n2617), .S0(n3055), .Y(prev_ReadData2[21]) );
  MX4X1 U639 ( .A(n2809), .B(n2807), .C(n2808), .D(n2806), .S0(n3059), .S1(
        n3064), .Y(n2617) );
  OAI2BB2XL U640 ( .B0(n3124), .B1(n3169), .A0N(prev_ReadData2[20]), .A1N(
        n3171), .Y(ReadData2[20]) );
  MXI2X1 U641 ( .A(n2614), .B(n2615), .S0(n3055), .Y(prev_ReadData2[20]) );
  MX4X1 U642 ( .A(n2801), .B(n2799), .C(n2800), .D(n2798), .S0(n3059), .S1(
        n3064), .Y(n2615) );
  OAI2BB2XL U643 ( .B0(n3112), .B1(n3169), .A0N(prev_ReadData2[26]), .A1N(
        n3170), .Y(ReadData2[26]) );
  MXI2X1 U644 ( .A(n2626), .B(n2627), .S0(n3055), .Y(prev_ReadData2[26]) );
  MX4X1 U645 ( .A(n2849), .B(n2847), .C(n2848), .D(n2846), .S0(n3060), .S1(
        n3061), .Y(n2627) );
  OAI2BB2XL U646 ( .B0(n3110), .B1(n3169), .A0N(prev_ReadData2[27]), .A1N(
        n3170), .Y(ReadData2[27]) );
  MXI2X1 U647 ( .A(n2628), .B(n2629), .S0(n3055), .Y(prev_ReadData2[27]) );
  MX4X1 U648 ( .A(n2857), .B(n2855), .C(n2856), .D(n2854), .S0(n3060), .S1(
        n3062), .Y(n2629) );
  OAI2BB2XL U649 ( .B0(n3114), .B1(n125), .A0N(prev_ReadData2[25]), .A1N(n3170), .Y(ReadData2[25]) );
  MXI2X1 U650 ( .A(n2624), .B(n2625), .S0(n3055), .Y(prev_ReadData2[25]) );
  MX4X1 U651 ( .A(n2841), .B(n2839), .C(n2840), .D(n2838), .S0(n3059), .S1(
        n3064), .Y(n2625) );
  OAI2BB2XL U652 ( .B0(n3116), .B1(n3170), .A0N(prev_ReadData2[24]), .A1N(
        n3171), .Y(ReadData2[24]) );
  MXI2X1 U653 ( .A(n2622), .B(n2623), .S0(n3055), .Y(prev_ReadData2[24]) );
  MX4X1 U654 ( .A(n2833), .B(n2831), .C(n2832), .D(n2830), .S0(n3059), .S1(
        n3064), .Y(n2623) );
  OAI2BB2XL U655 ( .B0(n3160), .B1(n125), .A0N(prev_ReadData2[2]), .A1N(n3171), 
        .Y(ReadData2[2]) );
  MXI2X1 U656 ( .A(n2578), .B(n2579), .S0(n3055), .Y(prev_ReadData2[2]) );
  MX4X1 U657 ( .A(n2661), .B(n2659), .C(n2660), .D(n2658), .S0(n3057), .S1(
        n3062), .Y(n2578) );
  OAI2BB2XL U658 ( .B0(n3162), .B1(n3169), .A0N(prev_ReadData2[1]), .A1N(n3171), .Y(ReadData2[1]) );
  MXI2X1 U659 ( .A(n2576), .B(n2577), .S0(n3055), .Y(prev_ReadData2[1]) );
  MX4X1 U660 ( .A(n2653), .B(n2651), .C(n2652), .D(n2650), .S0(n3060), .S1(
        n3061), .Y(n2576) );
  OAI2BB2XL U661 ( .B0(n3142), .B1(n3169), .A0N(prev_ReadData2[11]), .A1N(
        n3171), .Y(ReadData2[11]) );
  MXI2X1 U662 ( .A(n2596), .B(n2597), .S0(n3054), .Y(prev_ReadData2[11]) );
  MX4X1 U663 ( .A(n2733), .B(n2731), .C(n2732), .D(n2730), .S0(n3058), .S1(
        n3061), .Y(n2596) );
  OAI2BB2XL U664 ( .B0(n3144), .B1(n3169), .A0N(prev_ReadData2[10]), .A1N(
        n3171), .Y(ReadData2[10]) );
  MXI2X1 U665 ( .A(n2594), .B(n2595), .S0(n3054), .Y(prev_ReadData2[10]) );
  MX4X1 U666 ( .A(n2725), .B(n2723), .C(n2724), .D(n2722), .S0(n3058), .S1(
        n3061), .Y(n2594) );
  OAI2BB2XL U667 ( .B0(n3134), .B1(n3169), .A0N(prev_ReadData2[15]), .A1N(
        n3171), .Y(ReadData2[15]) );
  MXI2X1 U668 ( .A(n2604), .B(n2605), .S0(n3054), .Y(prev_ReadData2[15]) );
  MX4X1 U669 ( .A(n2765), .B(n2763), .C(n2764), .D(n2762), .S0(N10), .S1(n3063), .Y(n2604) );
  OAI2BB2XL U670 ( .B0(n3136), .B1(n3169), .A0N(prev_ReadData2[14]), .A1N(
        n3171), .Y(ReadData2[14]) );
  MXI2X1 U671 ( .A(n2602), .B(n2603), .S0(n3054), .Y(prev_ReadData2[14]) );
  MX4X1 U672 ( .A(n2757), .B(n2755), .C(n2756), .D(n2754), .S0(n3056), .S1(
        n3063), .Y(n2602) );
  OAI2BB2XL U673 ( .B0(n3138), .B1(n3169), .A0N(prev_ReadData2[13]), .A1N(
        n3169), .Y(ReadData2[13]) );
  MXI2X1 U674 ( .A(n2600), .B(n2601), .S0(n3054), .Y(prev_ReadData2[13]) );
  MX4X1 U675 ( .A(n2749), .B(n2747), .C(n2748), .D(n2746), .S0(n3058), .S1(
        n3061), .Y(n2600) );
  OAI2BB2XL U676 ( .B0(n3140), .B1(n3169), .A0N(prev_ReadData2[12]), .A1N(
        n3171), .Y(ReadData2[12]) );
  MXI2X1 U677 ( .A(n2598), .B(n2599), .S0(n3054), .Y(prev_ReadData2[12]) );
  MX4X1 U678 ( .A(n2741), .B(n2739), .C(n2740), .D(n2738), .S0(n3058), .S1(
        n3062), .Y(n2598) );
  OAI2BB2XL U679 ( .B0(n3116), .B1(n3167), .A0N(prev_ReadData1[24]), .A1N(
        n3168), .Y(ReadData1[24]) );
  MXI2X1 U680 ( .A(n63), .B(n65), .S0(n2527), .Y(prev_ReadData1[24]) );
  MX4X1 U681 ( .A(n2306), .B(n2304), .C(n2305), .D(n2303), .S0(n2532), .S1(
        n2536), .Y(n65) );
  OAI2BB2XL U682 ( .B0(n3124), .B1(n3166), .A0N(prev_ReadData1[20]), .A1N(
        n3168), .Y(ReadData1[20]) );
  MXI2X1 U683 ( .A(n42), .B(n46), .S0(n2527), .Y(prev_ReadData1[20]) );
  MX4X1 U684 ( .A(n2274), .B(n2272), .C(n2273), .D(n2271), .S0(n2532), .S1(
        n2536), .Y(n46) );
  OAI2BB2XL U685 ( .B0(n3132), .B1(n3166), .A0N(prev_ReadData1[16]), .A1N(
        n3168), .Y(ReadData1[16]) );
  MXI2X1 U686 ( .A(n34), .B(n35), .S0(n2528), .Y(prev_ReadData1[16]) );
  MX4X1 U687 ( .A(n2242), .B(n2240), .C(n2241), .D(n2239), .S0(n2531), .S1(
        n2535), .Y(n35) );
  OAI2BB2XL U688 ( .B0(n3140), .B1(n3166), .A0N(prev_ReadData1[12]), .A1N(
        n3168), .Y(ReadData1[12]) );
  MXI2X1 U689 ( .A(n26), .B(n27), .S0(N6), .Y(prev_ReadData1[12]) );
  MX4X1 U690 ( .A(n2214), .B(n2212), .C(n2213), .D(n2211), .S0(n2530), .S1(
        n2534), .Y(n26) );
  OAI2BB2XL U691 ( .B0(n3164), .B1(n3169), .A0N(prev_ReadData2[0]), .A1N(n3171), .Y(ReadData2[0]) );
  MXI2X1 U692 ( .A(n2574), .B(n2575), .S0(n3055), .Y(prev_ReadData2[0]) );
  MX4X1 U693 ( .A(n2641), .B(n2639), .C(n2640), .D(n2638), .S0(n3057), .S1(
        n3061), .Y(n2575) );
  CLKBUFX3 U694 ( .A(N6), .Y(n2528) );
  NOR2X2 U695 ( .A(n3443), .B(n3444), .Y(n58) );
  NOR2BX1 U696 ( .AN(n80), .B(n3441), .Y(n69) );
  NOR2BX1 U697 ( .AN(n100), .B(n3441), .Y(n89) );
  NOR2BX1 U698 ( .AN(n122), .B(n3441), .Y(n109) );
  NOR2BX1 U699 ( .AN(n59), .B(n3441), .Y(n44) );
  NOR2BX1 U700 ( .AN(n103), .B(n3442), .Y(n122) );
  CLKBUFX3 U701 ( .A(n9), .Y(n3292) );
  NAND2X1 U702 ( .A(n43), .B(n44), .Y(n9) );
  NAND2X1 U703 ( .A(n53), .B(n48), .Y(n51) );
  NAND2X1 U704 ( .A(n53), .B(n44), .Y(n54) );
  NAND2X1 U705 ( .A(n47), .B(n48), .Y(n45) );
  NAND2X1 U706 ( .A(n47), .B(n44), .Y(n49) );
  NAND2X1 U707 ( .A(n58), .B(n48), .Y(n56) );
  NAND2X1 U708 ( .A(n66), .B(n53), .Y(n74) );
  NAND2X1 U709 ( .A(n69), .B(n53), .Y(n76) );
  CLKBUFX3 U710 ( .A(n94), .Y(n3216) );
  NAND2X1 U711 ( .A(n86), .B(n53), .Y(n94) );
  NAND2X1 U712 ( .A(n89), .B(n53), .Y(n96) );
  NAND2X1 U713 ( .A(n106), .B(n53), .Y(n115) );
  NAND2X1 U714 ( .A(n109), .B(n53), .Y(n117) );
  NAND2X1 U715 ( .A(n66), .B(n47), .Y(n70) );
  NAND2X1 U716 ( .A(n69), .B(n47), .Y(n72) );
  NAND2X1 U717 ( .A(n66), .B(n58), .Y(n78) );
  NAND2X1 U718 ( .A(n86), .B(n47), .Y(n90) );
  NAND2X1 U719 ( .A(n89), .B(n47), .Y(n92) );
  NAND2X1 U720 ( .A(n86), .B(n58), .Y(n98) );
  NAND2X1 U721 ( .A(n106), .B(n47), .Y(n110) );
  NAND2X1 U722 ( .A(n109), .B(n47), .Y(n112) );
  NAND2X1 U723 ( .A(n106), .B(n58), .Y(n120) );
  NAND2X1 U724 ( .A(n66), .B(n43), .Y(n64) );
  NAND2X1 U725 ( .A(n86), .B(n43), .Y(n84) );
  NAND2X1 U726 ( .A(n106), .B(n43), .Y(n104) );
  NAND2X1 U727 ( .A(n69), .B(n43), .Y(n67) );
  NAND2X1 U728 ( .A(n89), .B(n43), .Y(n87) );
  NAND2X1 U729 ( .A(n109), .B(n43), .Y(n107) );
  MXI2X1 U730 ( .A(n1067), .B(n2367), .S0(n2570), .Y(n2370) );
  NOR2BX1 U731 ( .AN(n2548), .B(\register_r[3][31] ), .Y(n2367) );
  MX4X1 U732 ( .A(n2797), .B(n2795), .C(n2796), .D(n2794), .S0(n3056), .S1(
        n3063), .Y(n2612) );
  MXI4X1 U733 ( .A(\register_r[8][19] ), .B(\register_r[9][19] ), .C(
        \register_r[10][19] ), .D(\register_r[11][19] ), .S0(n3084), .S1(n3066), .Y(n2795) );
  MXI4X1 U734 ( .A(r_12[19]), .B(r_13[19]), .C(\register_r[14][19] ), .D(
        \register_r[15][19] ), .S0(n3084), .S1(n3066), .Y(n2794) );
  MXI4X1 U735 ( .A(\register_r[4][19] ), .B(\register_r[5][19] ), .C(
        \register_r[6][19] ), .D(\register_r[7][19] ), .S0(n3084), .S1(n3066), 
        .Y(n2796) );
  MX4X1 U736 ( .A(n2366), .B(n2364), .C(n2365), .D(n2363), .S0(n2533), .S1(
        n2537), .Y(n95) );
  MXI4X1 U737 ( .A(\register_r[8][31] ), .B(\register_r[9][31] ), .C(
        \register_r[10][31] ), .D(\register_r[11][31] ), .S0(n2557), .S1(n2540), .Y(n2364) );
  MXI4X1 U738 ( .A(r_12[31]), .B(r_13[31]), .C(\register_r[14][31] ), .D(
        \register_r[15][31] ), .S0(n2561), .S1(n2543), .Y(n2363) );
  NAND2X1 U739 ( .A(n2371), .B(n2370), .Y(n2366) );
  MX4X1 U740 ( .A(n2358), .B(n2356), .C(n2357), .D(n2355), .S0(n2533), .S1(
        n2537), .Y(n91) );
  MXI4X1 U741 ( .A(\register_r[8][30] ), .B(\register_r[9][30] ), .C(
        \register_r[10][30] ), .D(\register_r[11][30] ), .S0(n2560), .S1(n2542), .Y(n2356) );
  MXI4X1 U742 ( .A(r_12[30]), .B(r_13[30]), .C(\register_r[14][30] ), .D(
        \register_r[15][30] ), .S0(n2560), .S1(n2542), .Y(n2355) );
  MXI4X1 U743 ( .A(\register_r[4][30] ), .B(\register_r[5][30] ), .C(
        \register_r[6][30] ), .D(\register_r[7][30] ), .S0(n2561), .S1(n2542), 
        .Y(n2357) );
  MX4X1 U744 ( .A(n2350), .B(n2348), .C(n2349), .D(n2347), .S0(n2533), .S1(
        n2537), .Y(n85) );
  MXI4X1 U745 ( .A(\register_r[8][29] ), .B(\register_r[9][29] ), .C(
        \register_r[10][29] ), .D(\register_r[11][29] ), .S0(n2560), .S1(n2542), .Y(n2348) );
  MXI4X1 U746 ( .A(r_12[29]), .B(r_13[29]), .C(\register_r[14][29] ), .D(
        \register_r[15][29] ), .S0(n2560), .S1(n2542), .Y(n2347) );
  MXI4X1 U747 ( .A(\register_r[4][29] ), .B(\register_r[5][29] ), .C(
        \register_r[6][29] ), .D(\register_r[7][29] ), .S0(n2560), .S1(n2542), 
        .Y(n2349) );
  MX4X1 U748 ( .A(n2334), .B(n2332), .C(n2333), .D(n2331), .S0(n2533), .S1(
        n2537), .Y(n77) );
  MXI4X1 U749 ( .A(\register_r[8][27] ), .B(\register_r[9][27] ), .C(
        \register_r[10][27] ), .D(\register_r[11][27] ), .S0(n2559), .S1(n2541), .Y(n2332) );
  MXI4X1 U750 ( .A(r_12[27]), .B(r_13[27]), .C(\register_r[14][27] ), .D(
        \register_r[15][27] ), .S0(n2559), .S1(n2541), .Y(n2331) );
  MXI4X1 U751 ( .A(\register_r[4][27] ), .B(\register_r[5][27] ), .C(
        \register_r[6][27] ), .D(\register_r[7][27] ), .S0(n2559), .S1(n2541), 
        .Y(n2333) );
  MX4X1 U752 ( .A(n2326), .B(n2324), .C(n2325), .D(n2323), .S0(n2533), .S1(
        n2537), .Y(n73) );
  MXI4X1 U753 ( .A(\register_r[8][26] ), .B(\register_r[9][26] ), .C(
        \register_r[10][26] ), .D(\register_r[11][26] ), .S0(n2559), .S1(n2541), .Y(n2324) );
  MXI4X1 U754 ( .A(r_12[26]), .B(r_13[26]), .C(\register_r[14][26] ), .D(
        \register_r[15][26] ), .S0(n2559), .S1(n2541), .Y(n2323) );
  MXI4X1 U755 ( .A(\register_r[4][26] ), .B(\register_r[5][26] ), .C(
        \register_r[6][26] ), .D(\register_r[7][26] ), .S0(n2559), .S1(n2541), 
        .Y(n2325) );
  MX4X1 U756 ( .A(n2318), .B(n2316), .C(n2317), .D(n2315), .S0(n2532), .S1(
        n2536), .Y(n68) );
  MXI4X1 U757 ( .A(\register_r[8][25] ), .B(\register_r[9][25] ), .C(
        \register_r[10][25] ), .D(\register_r[11][25] ), .S0(n2558), .S1(n2541), .Y(n2316) );
  MXI4X1 U758 ( .A(r_12[25]), .B(r_13[25]), .C(\register_r[14][25] ), .D(
        \register_r[15][25] ), .S0(n2558), .S1(n2541), .Y(n2315) );
  MXI4X1 U759 ( .A(\register_r[4][25] ), .B(\register_r[5][25] ), .C(
        \register_r[6][25] ), .D(\register_r[7][25] ), .S0(n2558), .S1(n2541), 
        .Y(n2317) );
  MX4X1 U760 ( .A(n2302), .B(n2300), .C(n2301), .D(n2299), .S0(n2532), .S1(
        n2536), .Y(n61) );
  MXI4X1 U761 ( .A(\register_r[8][23] ), .B(\register_r[9][23] ), .C(
        \register_r[10][23] ), .D(\register_r[11][23] ), .S0(n2557), .S1(n2540), .Y(n2300) );
  MXI4X1 U762 ( .A(r_12[23]), .B(r_13[23]), .C(\register_r[14][23] ), .D(
        \register_r[15][23] ), .S0(n2557), .S1(n2540), .Y(n2299) );
  MXI4X1 U763 ( .A(\register_r[4][23] ), .B(\register_r[5][23] ), .C(
        \register_r[6][23] ), .D(\register_r[7][23] ), .S0(n2557), .S1(n2540), 
        .Y(n2301) );
  MX4X1 U764 ( .A(n2294), .B(n2292), .C(n2293), .D(n2291), .S0(n2532), .S1(
        n2536), .Y(n55) );
  MXI4X1 U765 ( .A(\register_r[8][22] ), .B(\register_r[9][22] ), .C(
        \register_r[10][22] ), .D(\register_r[11][22] ), .S0(n2557), .S1(n2540), .Y(n2292) );
  MXI4X1 U766 ( .A(r_12[22]), .B(r_13[22]), .C(\register_r[14][22] ), .D(
        \register_r[15][22] ), .S0(n2557), .S1(n2540), .Y(n2291) );
  MXI4X1 U767 ( .A(\register_r[4][22] ), .B(\register_r[5][22] ), .C(
        \register_r[6][22] ), .D(\register_r[7][22] ), .S0(n2557), .S1(n2540), 
        .Y(n2293) );
  MX4X1 U768 ( .A(n2286), .B(n2284), .C(n2285), .D(n2283), .S0(n2532), .S1(
        n2536), .Y(n50) );
  MXI4X1 U769 ( .A(\register_r[8][21] ), .B(\register_r[9][21] ), .C(
        \register_r[10][21] ), .D(\register_r[11][21] ), .S0(n2556), .S1(n2539), .Y(n2284) );
  MXI4X1 U770 ( .A(r_12[21]), .B(r_13[21]), .C(\register_r[14][21] ), .D(
        \register_r[15][21] ), .S0(n2556), .S1(n2539), .Y(n2283) );
  MXI4X1 U771 ( .A(\register_r[4][21] ), .B(\register_r[5][21] ), .C(
        \register_r[6][21] ), .D(\register_r[7][21] ), .S0(n2556), .S1(n2539), 
        .Y(n2285) );
  MX4X1 U772 ( .A(n2270), .B(n2268), .C(n2269), .D(n2267), .S0(n2531), .S1(
        n2535), .Y(n40) );
  MXI4X1 U773 ( .A(\register_r[8][19] ), .B(\register_r[9][19] ), .C(
        \register_r[10][19] ), .D(\register_r[11][19] ), .S0(n2555), .S1(n2539), .Y(n2268) );
  MXI4X1 U774 ( .A(r_12[19]), .B(r_13[19]), .C(\register_r[14][19] ), .D(
        \register_r[15][19] ), .S0(n2555), .S1(n2539), .Y(n2267) );
  MXI4X1 U775 ( .A(\register_r[4][19] ), .B(\register_r[5][19] ), .C(
        \register_r[6][19] ), .D(\register_r[7][19] ), .S0(n2555), .S1(n2539), 
        .Y(n2269) );
  MX4X1 U776 ( .A(n2262), .B(n2260), .C(n2261), .D(n2259), .S0(n2531), .S1(
        n2535), .Y(n38) );
  MXI4X1 U777 ( .A(\register_r[8][18] ), .B(\register_r[9][18] ), .C(
        \register_r[10][18] ), .D(\register_r[11][18] ), .S0(n2555), .S1(n2538), .Y(n2260) );
  MXI4X1 U778 ( .A(r_12[18]), .B(r_13[18]), .C(\register_r[14][18] ), .D(
        \register_r[15][18] ), .S0(n2555), .S1(n2538), .Y(n2259) );
  MXI4X1 U779 ( .A(\register_r[4][18] ), .B(\register_r[5][18] ), .C(
        \register_r[6][18] ), .D(\register_r[7][18] ), .S0(n2555), .S1(n2538), 
        .Y(n2261) );
  MX4X1 U780 ( .A(n2254), .B(n2252), .C(n2253), .D(n2251), .S0(n2531), .S1(
        n2535), .Y(n36) );
  MXI4X1 U781 ( .A(\register_r[8][17] ), .B(\register_r[9][17] ), .C(
        \register_r[10][17] ), .D(\register_r[11][17] ), .S0(n2554), .S1(n2538), .Y(n2252) );
  MXI4X1 U782 ( .A(r_12[17]), .B(r_13[17]), .C(\register_r[14][17] ), .D(
        \register_r[15][17] ), .S0(n2554), .S1(n2538), .Y(n2251) );
  MXI4X1 U783 ( .A(\register_r[4][17] ), .B(\register_r[5][17] ), .C(
        \register_r[6][17] ), .D(\register_r[7][17] ), .S0(n2554), .S1(n2538), 
        .Y(n2253) );
  MX4X1 U784 ( .A(n116), .B(n113), .C(n114), .D(n111), .S0(n2530), .S1(n2537), 
        .Y(n1) );
  MXI4X1 U785 ( .A(\register_r[8][0] ), .B(\register_r[9][0] ), .C(
        \register_r[10][0] ), .D(\register_r[11][0] ), .S0(n2561), .S1(n2543), 
        .Y(n113) );
  MXI4X1 U786 ( .A(r_12[0]), .B(r_13[0]), .C(\register_r[14][0] ), .D(
        \register_r[15][0] ), .S0(n2561), .S1(n2543), .Y(n111) );
  MXI4X1 U787 ( .A(\register_r[4][0] ), .B(\register_r[5][0] ), .C(
        \register_r[6][0] ), .D(\register_r[7][0] ), .S0(n2561), .S1(n2543), 
        .Y(n114) );
  MX4X1 U788 ( .A(n2234), .B(n2232), .C(n2233), .D(n2231), .S0(n2531), .S1(
        n2535), .Y(n33) );
  MXI4X1 U789 ( .A(\register_r[16][15] ), .B(\register_r[17][15] ), .C(
        \register_r[18][15] ), .D(\register_r[19][15] ), .S0(n2568), .S1(n2546), .Y(n2234) );
  MXI4X1 U790 ( .A(\register_r[24][15] ), .B(\register_r[25][15] ), .C(
        \register_r[26][15] ), .D(\register_r[27][15] ), .S0(n2568), .S1(n2546), .Y(n2232) );
  MXI4X1 U791 ( .A(\register_r[28][15] ), .B(\register_r[29][15] ), .C(
        \register_r[30][15] ), .D(\register_r[31][15] ), .S0(n2568), .S1(n2546), .Y(n2231) );
  MX4X1 U792 ( .A(n2226), .B(n2224), .C(n2225), .D(n2223), .S0(n2531), .S1(
        n2535), .Y(n31) );
  MXI4X1 U793 ( .A(\register_r[16][14] ), .B(\register_r[17][14] ), .C(
        \register_r[18][14] ), .D(\register_r[19][14] ), .S0(n2568), .S1(n2546), .Y(n2226) );
  MXI4X1 U794 ( .A(\register_r[24][14] ), .B(\register_r[25][14] ), .C(
        \register_r[26][14] ), .D(\register_r[27][14] ), .S0(n2568), .S1(n2546), .Y(n2224) );
  MXI4X1 U795 ( .A(\register_r[28][14] ), .B(\register_r[29][14] ), .C(
        \register_r[30][14] ), .D(\register_r[31][14] ), .S0(n2567), .S1(n2546), .Y(n2223) );
  MX4X1 U796 ( .A(n2218), .B(n2216), .C(n2217), .D(n2215), .S0(n2530), .S1(
        n2534), .Y(n29) );
  MXI4X1 U797 ( .A(\register_r[16][13] ), .B(\register_r[17][13] ), .C(
        \register_r[18][13] ), .D(\register_r[19][13] ), .S0(n2567), .S1(n2546), .Y(n2218) );
  MXI4X1 U798 ( .A(\register_r[24][13] ), .B(\register_r[25][13] ), .C(
        \register_r[26][13] ), .D(\register_r[27][13] ), .S0(n2567), .S1(n2546), .Y(n2216) );
  MXI4X1 U799 ( .A(\register_r[28][13] ), .B(\register_r[29][13] ), .C(
        \register_r[30][13] ), .D(\register_r[31][13] ), .S0(n2567), .S1(n2546), .Y(n2215) );
  MX4X1 U800 ( .A(n2202), .B(n2200), .C(n2201), .D(n2199), .S0(n2530), .S1(
        n2536), .Y(n25) );
  MXI4X1 U801 ( .A(\register_r[16][11] ), .B(\register_r[17][11] ), .C(
        \register_r[18][11] ), .D(\register_r[19][11] ), .S0(n2566), .S1(n2545), .Y(n2202) );
  MXI4X1 U802 ( .A(\register_r[24][11] ), .B(\register_r[25][11] ), .C(
        \register_r[26][11] ), .D(\register_r[27][11] ), .S0(n2566), .S1(n2545), .Y(n2200) );
  MXI4X1 U803 ( .A(\register_r[28][11] ), .B(\register_r[29][11] ), .C(
        \register_r[30][11] ), .D(\register_r[31][11] ), .S0(n2566), .S1(n2545), .Y(n2199) );
  MX4X1 U804 ( .A(n2194), .B(n2192), .C(n2193), .D(n2191), .S0(n2530), .S1(
        n2535), .Y(n23) );
  MXI4X1 U805 ( .A(\register_r[16][10] ), .B(\register_r[17][10] ), .C(
        \register_r[18][10] ), .D(\register_r[19][10] ), .S0(n2566), .S1(n2545), .Y(n2194) );
  MXI4X1 U806 ( .A(\register_r[24][10] ), .B(\register_r[25][10] ), .C(
        \register_r[26][10] ), .D(\register_r[27][10] ), .S0(n2566), .S1(n2545), .Y(n2192) );
  MXI4X1 U807 ( .A(\register_r[28][10] ), .B(\register_r[29][10] ), .C(
        \register_r[30][10] ), .D(\register_r[31][10] ), .S0(n2566), .S1(n2545), .Y(n2191) );
  MX4X1 U808 ( .A(n2186), .B(n2184), .C(n2185), .D(n2183), .S0(n2530), .S1(
        n2534), .Y(n21) );
  MXI4X1 U809 ( .A(\register_r[16][9] ), .B(\register_r[17][9] ), .C(
        \register_r[18][9] ), .D(\register_r[19][9] ), .S0(n2565), .S1(n2545), 
        .Y(n2186) );
  MXI4X1 U810 ( .A(\register_r[24][9] ), .B(\register_r[25][9] ), .C(
        \register_r[26][9] ), .D(\register_r[27][9] ), .S0(n2565), .S1(n2545), 
        .Y(n2184) );
  MXI4X1 U811 ( .A(\register_r[28][9] ), .B(\register_r[29][9] ), .C(
        \register_r[30][9] ), .D(\register_r[31][9] ), .S0(n2565), .S1(n2544), 
        .Y(n2183) );
  MX4X1 U812 ( .A(n2170), .B(n2168), .C(n2169), .D(n2167), .S0(n2533), .S1(
        n2534), .Y(n17) );
  MXI4X1 U813 ( .A(\register_r[16][7] ), .B(\register_r[17][7] ), .C(
        \register_r[18][7] ), .D(\register_r[19][7] ), .S0(n2564), .S1(n2544), 
        .Y(n2170) );
  MXI4X1 U814 ( .A(\register_r[24][7] ), .B(\register_r[25][7] ), .C(
        \register_r[26][7] ), .D(\register_r[27][7] ), .S0(n2564), .S1(n2544), 
        .Y(n2168) );
  MXI4X1 U815 ( .A(\register_r[28][7] ), .B(\register_r[29][7] ), .C(
        \register_r[30][7] ), .D(\register_r[31][7] ), .S0(n2564), .S1(n2544), 
        .Y(n2167) );
  MX4X1 U816 ( .A(n2162), .B(n2160), .C(n2161), .D(n2159), .S0(n2529), .S1(
        n2534), .Y(n15) );
  MXI4X1 U817 ( .A(\register_r[16][6] ), .B(\register_r[17][6] ), .C(
        \register_r[18][6] ), .D(\register_r[19][6] ), .S0(n2564), .S1(n2544), 
        .Y(n2162) );
  MXI4X1 U818 ( .A(\register_r[24][6] ), .B(\register_r[25][6] ), .C(
        \register_r[26][6] ), .D(\register_r[27][6] ), .S0(n2564), .S1(n2544), 
        .Y(n2160) );
  MXI4X1 U819 ( .A(\register_r[28][6] ), .B(\register_r[29][6] ), .C(
        \register_r[30][6] ), .D(\register_r[31][6] ), .S0(n2564), .S1(n2541), 
        .Y(n2159) );
  MX4X1 U820 ( .A(n2154), .B(n2152), .C(n2153), .D(n2151), .S0(n2529), .S1(
        n2536), .Y(n13) );
  MXI4X1 U821 ( .A(\register_r[16][5] ), .B(\register_r[17][5] ), .C(
        \register_r[18][5] ), .D(\register_r[19][5] ), .S0(n2563), .S1(n2551), 
        .Y(n2154) );
  MXI4X1 U822 ( .A(\register_r[24][5] ), .B(\register_r[25][5] ), .C(
        \register_r[26][5] ), .D(\register_r[27][5] ), .S0(n2563), .S1(N3), 
        .Y(n2152) );
  MXI4X1 U823 ( .A(\register_r[28][5] ), .B(\register_r[29][5] ), .C(
        \register_r[30][5] ), .D(\register_r[31][5] ), .S0(n2563), .S1(n2551), 
        .Y(n2151) );
  MX4X1 U824 ( .A(n2138), .B(n2136), .C(n2137), .D(n2135), .S0(n2529), .S1(
        n2534), .Y(n8) );
  MXI4X1 U825 ( .A(\register_r[16][3] ), .B(\register_r[17][3] ), .C(
        \register_r[18][3] ), .D(\register_r[19][3] ), .S0(n2563), .S1(n2550), 
        .Y(n2138) );
  MXI4X1 U826 ( .A(\register_r[24][3] ), .B(\register_r[25][3] ), .C(
        \register_r[26][3] ), .D(\register_r[27][3] ), .S0(n2562), .S1(n2544), 
        .Y(n2136) );
  MXI4X1 U827 ( .A(\register_r[28][3] ), .B(\register_r[29][3] ), .C(
        \register_r[30][3] ), .D(\register_r[31][3] ), .S0(n2562), .S1(n2546), 
        .Y(n2135) );
  MX4X1 U828 ( .A(n2130), .B(n2128), .C(n2129), .D(n2127), .S0(n2529), .S1(
        n2535), .Y(n6) );
  MXI4X1 U829 ( .A(\register_r[16][2] ), .B(\register_r[17][2] ), .C(
        \register_r[18][2] ), .D(\register_r[19][2] ), .S0(n2562), .S1(n2543), 
        .Y(n2130) );
  MXI4X1 U830 ( .A(\register_r[24][2] ), .B(\register_r[25][2] ), .C(
        \register_r[26][2] ), .D(\register_r[27][2] ), .S0(n2562), .S1(n2543), 
        .Y(n2128) );
  MXI4X1 U831 ( .A(\register_r[28][2] ), .B(\register_r[29][2] ), .C(
        \register_r[30][2] ), .D(\register_r[31][2] ), .S0(n2562), .S1(n2543), 
        .Y(n2127) );
  MX4X1 U832 ( .A(n124), .B(n119), .C(n121), .D(n118), .S0(n2529), .S1(n2535), 
        .Y(n4) );
  MXI4X1 U833 ( .A(\register_r[24][1] ), .B(\register_r[25][1] ), .C(
        \register_r[26][1] ), .D(\register_r[27][1] ), .S0(n2561), .S1(n2543), 
        .Y(n119) );
  MXI4X1 U834 ( .A(\register_r[16][1] ), .B(\register_r[17][1] ), .C(
        \register_r[18][1] ), .D(\register_r[19][1] ), .S0(n2562), .S1(n2543), 
        .Y(n124) );
  MXI4X1 U835 ( .A(\register_r[28][1] ), .B(\register_r[29][1] ), .C(
        \register_r[30][1] ), .D(\register_r[31][1] ), .S0(n2561), .S1(n2543), 
        .Y(n118) );
  NOR2BX1 U836 ( .AN(n3074), .B(\register_r[3][19] ), .Y(n2954) );
  NOR2BX1 U837 ( .AN(n2548), .B(\register_r[3][30] ), .Y(n2372) );
  NOR2BX1 U838 ( .AN(n2548), .B(\register_r[3][29] ), .Y(n2377) );
  NOR2BX1 U839 ( .AN(n2548), .B(\register_r[3][27] ), .Y(n2387) );
  NOR2BX1 U840 ( .AN(n2548), .B(\register_r[3][26] ), .Y(n2392) );
  NOR2BX1 U841 ( .AN(n2548), .B(\register_r[3][25] ), .Y(n2397) );
  NOR2BX1 U842 ( .AN(n2547), .B(\register_r[3][23] ), .Y(n2407) );
  NOR2BX1 U843 ( .AN(n2547), .B(\register_r[3][22] ), .Y(n2412) );
  NOR2BX1 U844 ( .AN(n2547), .B(\register_r[3][21] ), .Y(n2417) );
  NOR2BX1 U845 ( .AN(n2547), .B(\register_r[3][19] ), .Y(n2427) );
  NOR2BX1 U846 ( .AN(n2547), .B(\register_r[3][18] ), .Y(n2432) );
  NOR2BX1 U847 ( .AN(n2547), .B(\register_r[3][17] ), .Y(n2437) );
  NOR2BX1 U848 ( .AN(n2547), .B(\register_r[3][15] ), .Y(n2447) );
  NOR2BX1 U849 ( .AN(n2547), .B(\register_r[3][14] ), .Y(n2452) );
  NOR2BX1 U850 ( .AN(n2547), .B(\register_r[3][13] ), .Y(n2457) );
  NOR2BX1 U851 ( .AN(n2547), .B(\register_r[3][11] ), .Y(n2467) );
  NOR2BX1 U852 ( .AN(n2547), .B(\register_r[3][10] ), .Y(n2472) );
  NOR2BX1 U853 ( .AN(n2547), .B(\register_r[3][9] ), .Y(n2477) );
  NOR2BX1 U854 ( .AN(n2547), .B(\register_r[3][7] ), .Y(n2487) );
  NOR2BX1 U855 ( .AN(n2548), .B(\register_r[3][6] ), .Y(n2492) );
  NOR2BX1 U856 ( .AN(n2547), .B(\register_r[3][5] ), .Y(n2497) );
  NOR2BX1 U857 ( .AN(n2548), .B(\register_r[3][3] ), .Y(n2507) );
  NOR2BX1 U858 ( .AN(n2548), .B(\register_r[3][2] ), .Y(n2512) );
  NOR2BX1 U859 ( .AN(n2548), .B(\register_r[3][1] ), .Y(n2517) );
  NOR2BX1 U860 ( .AN(n2548), .B(\register_r[3][0] ), .Y(n2522) );
  NAND2X1 U861 ( .A(n2521), .B(n2520), .Y(n2126) );
  NOR2X1 U862 ( .A(n2519), .B(n2518), .Y(n2521) );
  MXI2X1 U863 ( .A(n1097), .B(n2517), .S0(n2568), .Y(n2520) );
  NOR2X1 U864 ( .A(n2550), .B(\register_r[1][1] ), .Y(n2519) );
  NAND2X1 U865 ( .A(n2958), .B(n2957), .Y(n2797) );
  NOR2X1 U866 ( .A(n2956), .B(n2955), .Y(n2958) );
  MXI2X1 U867 ( .A(n1079), .B(n2954), .S0(n3098), .Y(n2957) );
  NOR2X1 U868 ( .A(n3079), .B(\register_r[1][19] ), .Y(n2956) );
  NAND2X1 U869 ( .A(n2381), .B(n2380), .Y(n2350) );
  NOR2X1 U870 ( .A(n2379), .B(n2378), .Y(n2381) );
  MXI2X1 U871 ( .A(n1069), .B(n2377), .S0(n2570), .Y(n2380) );
  NOR2X1 U872 ( .A(n2543), .B(\register_r[1][29] ), .Y(n2379) );
  NAND2X1 U873 ( .A(n2396), .B(n2395), .Y(n2326) );
  NOR2X1 U874 ( .A(n2394), .B(n2393), .Y(n2396) );
  MXI2X1 U875 ( .A(n1072), .B(n2392), .S0(n2570), .Y(n2395) );
  NOR2X1 U876 ( .A(n2550), .B(n2572), .Y(n2393) );
  NAND2X1 U877 ( .A(n2411), .B(n2410), .Y(n2302) );
  NOR2X1 U878 ( .A(n2409), .B(n2408), .Y(n2411) );
  MXI2X1 U879 ( .A(n1075), .B(n2407), .S0(n2570), .Y(n2410) );
  NOR2X1 U880 ( .A(n2549), .B(\register_r[1][23] ), .Y(n2409) );
  NAND2X1 U881 ( .A(n2416), .B(n2415), .Y(n2294) );
  NOR2X1 U882 ( .A(n2414), .B(n2413), .Y(n2416) );
  MXI2X1 U883 ( .A(n1076), .B(n2412), .S0(n2570), .Y(n2415) );
  NOR2X1 U884 ( .A(n2549), .B(\register_r[1][22] ), .Y(n2414) );
  NAND2X1 U885 ( .A(n2421), .B(n2420), .Y(n2286) );
  NOR2X1 U886 ( .A(n2419), .B(n2418), .Y(n2421) );
  MXI2X1 U887 ( .A(n1077), .B(n2417), .S0(n2570), .Y(n2420) );
  NOR2X1 U888 ( .A(n2540), .B(\register_r[1][21] ), .Y(n2419) );
  NAND2X1 U889 ( .A(n2431), .B(n2430), .Y(n2270) );
  NOR2X1 U890 ( .A(n2429), .B(n2428), .Y(n2431) );
  MXI2X1 U891 ( .A(n1079), .B(n2427), .S0(n2570), .Y(n2430) );
  NOR2X1 U892 ( .A(n2545), .B(\register_r[1][19] ), .Y(n2429) );
  NAND2X1 U893 ( .A(n2436), .B(n2435), .Y(n2262) );
  NOR2X1 U894 ( .A(n2434), .B(n2433), .Y(n2436) );
  MXI2X1 U895 ( .A(n1080), .B(n2432), .S0(n2570), .Y(n2435) );
  NOR2X1 U896 ( .A(n2540), .B(\register_r[1][18] ), .Y(n2434) );
  NAND2X1 U897 ( .A(n2441), .B(n2440), .Y(n2254) );
  NOR2X1 U898 ( .A(n2439), .B(n2438), .Y(n2441) );
  MXI2X1 U899 ( .A(n1081), .B(n2437), .S0(n2570), .Y(n2440) );
  NOR2X1 U900 ( .A(n2546), .B(\register_r[1][17] ), .Y(n2439) );
  NAND2X1 U901 ( .A(n2451), .B(n2450), .Y(n2238) );
  NOR2X1 U902 ( .A(n2449), .B(n2448), .Y(n2451) );
  MXI2X1 U903 ( .A(n1083), .B(n2447), .S0(n2570), .Y(n2450) );
  NOR2X1 U904 ( .A(n2546), .B(\register_r[1][15] ), .Y(n2449) );
  NAND2X1 U905 ( .A(n2456), .B(n2455), .Y(n2230) );
  NOR2X1 U906 ( .A(n2454), .B(n2453), .Y(n2456) );
  MXI2X1 U907 ( .A(n1084), .B(n2452), .S0(n2569), .Y(n2455) );
  NOR2X1 U908 ( .A(n2550), .B(\register_r[1][14] ), .Y(n2454) );
  NAND2X1 U909 ( .A(n2461), .B(n2460), .Y(n2222) );
  NOR2X1 U910 ( .A(n2459), .B(n2458), .Y(n2461) );
  MXI2X1 U911 ( .A(n1085), .B(n2457), .S0(n2569), .Y(n2460) );
  NOR2X1 U912 ( .A(n2550), .B(\register_r[1][13] ), .Y(n2459) );
  NAND2X1 U913 ( .A(n2471), .B(n2470), .Y(n2206) );
  NOR2X1 U914 ( .A(n2469), .B(n2468), .Y(n2471) );
  MXI2X1 U915 ( .A(n1087), .B(n2467), .S0(n2569), .Y(n2470) );
  NOR2X1 U916 ( .A(n2550), .B(\register_r[1][11] ), .Y(n2469) );
  NAND2X1 U917 ( .A(n2476), .B(n2475), .Y(n2198) );
  NOR2X1 U918 ( .A(n2474), .B(n2473), .Y(n2476) );
  MXI2X1 U919 ( .A(n1088), .B(n2472), .S0(n2569), .Y(n2475) );
  NOR2X1 U920 ( .A(n2549), .B(\register_r[1][10] ), .Y(n2474) );
  NAND2X1 U921 ( .A(n2481), .B(n2480), .Y(n2190) );
  NOR2X1 U922 ( .A(n2479), .B(n2478), .Y(n2481) );
  MXI2X1 U923 ( .A(n1089), .B(n2477), .S0(n2569), .Y(n2480) );
  NOR2X1 U924 ( .A(n2549), .B(\register_r[1][9] ), .Y(n2479) );
  NAND2X1 U925 ( .A(n2491), .B(n2490), .Y(n2174) );
  NOR2X1 U926 ( .A(n2489), .B(n2488), .Y(n2491) );
  MXI2X1 U927 ( .A(n1091), .B(n2487), .S0(n2569), .Y(n2490) );
  NOR2X1 U928 ( .A(n2549), .B(\register_r[1][7] ), .Y(n2489) );
  NAND2X1 U929 ( .A(n2496), .B(n2495), .Y(n2166) );
  NOR2X1 U930 ( .A(n2494), .B(n2493), .Y(n2496) );
  MXI2X1 U931 ( .A(n1092), .B(n2492), .S0(n2569), .Y(n2495) );
  NOR2X1 U932 ( .A(n2548), .B(\register_r[1][6] ), .Y(n2494) );
  NAND2X1 U933 ( .A(n2501), .B(n2500), .Y(n2158) );
  NOR2X1 U934 ( .A(n2499), .B(n2498), .Y(n2501) );
  MXI2X1 U935 ( .A(n1093), .B(n2497), .S0(n2569), .Y(n2500) );
  NOR2X1 U936 ( .A(n2549), .B(\register_r[1][5] ), .Y(n2499) );
  NAND2X1 U937 ( .A(n2511), .B(n2510), .Y(n2142) );
  NOR2X1 U938 ( .A(n2509), .B(n2508), .Y(n2511) );
  MXI2X1 U939 ( .A(n1095), .B(n2507), .S0(n2569), .Y(n2510) );
  NOR2X1 U940 ( .A(n2549), .B(\register_r[1][3] ), .Y(n2509) );
  NAND2X1 U941 ( .A(n2516), .B(n2515), .Y(n2134) );
  NOR2X1 U942 ( .A(n2514), .B(n2513), .Y(n2516) );
  MXI2X1 U943 ( .A(n1096), .B(n2512), .S0(n2569), .Y(n2515) );
  NOR2X1 U944 ( .A(n2550), .B(\register_r[1][2] ), .Y(n2514) );
  NAND2X1 U945 ( .A(n2376), .B(n2375), .Y(n2358) );
  NOR2X1 U946 ( .A(n2374), .B(n2373), .Y(n2376) );
  MXI2X1 U947 ( .A(n1068), .B(n2372), .S0(n2571), .Y(n2375) );
  NOR2X1 U948 ( .A(n2550), .B(\register_r[1][30] ), .Y(n2374) );
  NAND2X1 U949 ( .A(n2391), .B(n2390), .Y(n2334) );
  NOR2X1 U950 ( .A(n2389), .B(n2388), .Y(n2391) );
  MXI2X1 U951 ( .A(n1071), .B(n2387), .S0(n2571), .Y(n2390) );
  NOR2X1 U952 ( .A(n2550), .B(\register_r[1][27] ), .Y(n2389) );
  NAND2X1 U953 ( .A(n2401), .B(n2400), .Y(n2318) );
  NOR2X1 U954 ( .A(n2399), .B(n2398), .Y(n2401) );
  MXI2X1 U955 ( .A(n1073), .B(n2397), .S0(n2571), .Y(n2400) );
  NOR2X1 U956 ( .A(n2546), .B(\register_r[1][25] ), .Y(n2399) );
  NAND2X1 U957 ( .A(n2526), .B(n2525), .Y(n116) );
  NOR2X1 U958 ( .A(n2524), .B(n2523), .Y(n2526) );
  MXI2X1 U959 ( .A(n1098), .B(n2522), .S0(n2571), .Y(n2525) );
  NOR2X1 U960 ( .A(n2543), .B(\register_r[1][0] ), .Y(n2524) );
  MXI4X1 U961 ( .A(\register_r[4][31] ), .B(\register_r[5][31] ), .C(
        \register_r[6][31] ), .D(\register_r[7][31] ), .S0(n2568), .S1(n2547), 
        .Y(n2365) );
  MXI4X1 U962 ( .A(\register_r[20][31] ), .B(\register_r[21][31] ), .C(
        \register_r[22][31] ), .D(\register_r[23][31] ), .S0(n2561), .S1(n2542), .Y(n2361) );
  MXI4X1 U963 ( .A(\register_r[20][30] ), .B(\register_r[21][30] ), .C(
        \register_r[22][30] ), .D(\register_r[23][30] ), .S0(n2560), .S1(n2542), .Y(n2353) );
  MXI4X1 U964 ( .A(\register_r[20][29] ), .B(\register_r[21][29] ), .C(
        \register_r[22][29] ), .D(\register_r[23][29] ), .S0(n2560), .S1(n2542), .Y(n2345) );
  MXI4X1 U965 ( .A(\register_r[20][27] ), .B(\register_r[21][27] ), .C(
        \register_r[22][27] ), .D(\register_r[23][27] ), .S0(n2559), .S1(n2541), .Y(n2329) );
  MXI4X1 U966 ( .A(\register_r[20][26] ), .B(\register_r[21][26] ), .C(
        \register_r[22][26] ), .D(\register_r[23][26] ), .S0(n2558), .S1(n2541), .Y(n2321) );
  MXI4X1 U967 ( .A(\register_r[20][25] ), .B(\register_r[21][25] ), .C(
        \register_r[22][25] ), .D(\register_r[23][25] ), .S0(n2558), .S1(n2541), .Y(n2313) );
  MXI4X1 U968 ( .A(\register_r[20][23] ), .B(\register_r[21][23] ), .C(
        \register_r[22][23] ), .D(\register_r[23][23] ), .S0(n2557), .S1(n2540), .Y(n2297) );
  MXI4X1 U969 ( .A(\register_r[20][22] ), .B(\register_r[21][22] ), .C(
        \register_r[22][22] ), .D(\register_r[23][22] ), .S0(n2556), .S1(n2540), .Y(n2289) );
  MXI4X1 U970 ( .A(\register_r[20][21] ), .B(\register_r[21][21] ), .C(
        \register_r[22][21] ), .D(\register_r[23][21] ), .S0(n2556), .S1(n2539), .Y(n2281) );
  MXI4X1 U971 ( .A(\register_r[20][19] ), .B(\register_r[21][19] ), .C(
        \register_r[22][19] ), .D(\register_r[23][19] ), .S0(n2555), .S1(n2539), .Y(n2265) );
  MXI4X1 U972 ( .A(\register_r[20][18] ), .B(\register_r[21][18] ), .C(
        \register_r[22][18] ), .D(\register_r[23][18] ), .S0(n2555), .S1(n2538), .Y(n2257) );
  MXI4X1 U973 ( .A(\register_r[20][17] ), .B(\register_r[21][17] ), .C(
        \register_r[22][17] ), .D(\register_r[23][17] ), .S0(n2554), .S1(n2538), .Y(n2249) );
  MXI4X1 U974 ( .A(\register_r[20][15] ), .B(\register_r[21][15] ), .C(
        \register_r[22][15] ), .D(\register_r[23][15] ), .S0(n2568), .S1(n2546), .Y(n2233) );
  MXI4X1 U975 ( .A(\register_r[4][15] ), .B(\register_r[5][15] ), .C(
        \register_r[6][15] ), .D(\register_r[7][15] ), .S0(n2565), .S1(n2544), 
        .Y(n2237) );
  MXI4X1 U976 ( .A(\register_r[20][14] ), .B(\register_r[21][14] ), .C(
        \register_r[22][14] ), .D(\register_r[23][14] ), .S0(n2568), .S1(n2546), .Y(n2225) );
  MXI4X1 U977 ( .A(\register_r[4][14] ), .B(\register_r[5][14] ), .C(
        \register_r[6][14] ), .D(\register_r[7][14] ), .S0(n2568), .S1(n2546), 
        .Y(n2229) );
  MXI4X1 U978 ( .A(\register_r[20][13] ), .B(\register_r[21][13] ), .C(
        \register_r[22][13] ), .D(\register_r[23][13] ), .S0(n2567), .S1(n2546), .Y(n2217) );
  MXI4X1 U979 ( .A(\register_r[4][13] ), .B(\register_r[5][13] ), .C(
        \register_r[6][13] ), .D(\register_r[7][13] ), .S0(n2567), .S1(n2546), 
        .Y(n2221) );
  MXI4X1 U980 ( .A(\register_r[20][11] ), .B(\register_r[21][11] ), .C(
        \register_r[22][11] ), .D(\register_r[23][11] ), .S0(n2566), .S1(n2545), .Y(n2201) );
  MXI4X1 U981 ( .A(\register_r[4][11] ), .B(\register_r[5][11] ), .C(
        \register_r[6][11] ), .D(\register_r[7][11] ), .S0(n2567), .S1(n2545), 
        .Y(n2205) );
  MXI4X1 U982 ( .A(\register_r[20][10] ), .B(\register_r[21][10] ), .C(
        \register_r[22][10] ), .D(\register_r[23][10] ), .S0(n2566), .S1(n2545), .Y(n2193) );
  MXI4X1 U983 ( .A(\register_r[4][10] ), .B(\register_r[5][10] ), .C(
        \register_r[6][10] ), .D(\register_r[7][10] ), .S0(n2566), .S1(n2545), 
        .Y(n2197) );
  MXI4X1 U984 ( .A(\register_r[20][9] ), .B(\register_r[21][9] ), .C(
        \register_r[22][9] ), .D(\register_r[23][9] ), .S0(n2565), .S1(n2545), 
        .Y(n2185) );
  MXI4X1 U985 ( .A(\register_r[4][9] ), .B(\register_r[5][9] ), .C(
        \register_r[6][9] ), .D(\register_r[7][9] ), .S0(n2566), .S1(n2545), 
        .Y(n2189) );
  MXI4X1 U986 ( .A(\register_r[20][7] ), .B(\register_r[21][7] ), .C(
        \register_r[22][7] ), .D(\register_r[23][7] ), .S0(n2564), .S1(n2544), 
        .Y(n2169) );
  MXI4X1 U987 ( .A(\register_r[4][7] ), .B(\register_r[5][7] ), .C(
        \register_r[6][7] ), .D(\register_r[7][7] ), .S0(n2565), .S1(n2544), 
        .Y(n2173) );
  MXI4X1 U988 ( .A(\register_r[20][6] ), .B(\register_r[21][6] ), .C(
        \register_r[22][6] ), .D(\register_r[23][6] ), .S0(n2564), .S1(n2544), 
        .Y(n2161) );
  MXI4X1 U989 ( .A(\register_r[4][6] ), .B(\register_r[5][6] ), .C(
        \register_r[6][6] ), .D(\register_r[7][6] ), .S0(n2564), .S1(n2544), 
        .Y(n2165) );
  MXI4X1 U990 ( .A(\register_r[20][5] ), .B(\register_r[21][5] ), .C(
        \register_r[22][5] ), .D(\register_r[23][5] ), .S0(n2563), .S1(n2551), 
        .Y(n2153) );
  MXI4X1 U991 ( .A(\register_r[4][5] ), .B(\register_r[5][5] ), .C(
        \register_r[6][5] ), .D(\register_r[7][5] ), .S0(n2564), .S1(n2551), 
        .Y(n2157) );
  MXI4X1 U992 ( .A(\register_r[20][3] ), .B(\register_r[21][3] ), .C(
        \register_r[22][3] ), .D(\register_r[23][3] ), .S0(n2562), .S1(n2542), 
        .Y(n2137) );
  MXI4X1 U993 ( .A(\register_r[4][3] ), .B(\register_r[5][3] ), .C(
        \register_r[6][3] ), .D(\register_r[7][3] ), .S0(n2563), .S1(n2550), 
        .Y(n2141) );
  MXI4X1 U994 ( .A(\register_r[20][2] ), .B(\register_r[21][2] ), .C(
        \register_r[22][2] ), .D(\register_r[23][2] ), .S0(n2562), .S1(n2543), 
        .Y(n2129) );
  MXI4X1 U995 ( .A(\register_r[4][2] ), .B(\register_r[5][2] ), .C(
        \register_r[6][2] ), .D(\register_r[7][2] ), .S0(n2562), .S1(n2543), 
        .Y(n2133) );
  MXI4X1 U996 ( .A(\register_r[20][1] ), .B(\register_r[21][1] ), .C(
        \register_r[22][1] ), .D(\register_r[23][1] ), .S0(n2562), .S1(n2543), 
        .Y(n121) );
  MXI4X1 U997 ( .A(\register_r[4][1] ), .B(\register_r[5][1] ), .C(
        \register_r[6][1] ), .D(\register_r[7][1] ), .S0(n2562), .S1(n2543), 
        .Y(n2125) );
  MXI4X1 U998 ( .A(\register_r[20][0] ), .B(\register_r[21][0] ), .C(
        \register_r[22][0] ), .D(\register_r[23][0] ), .S0(n2561), .S1(n2543), 
        .Y(n105) );
  MXI4X1 U999 ( .A(\register_r[16][31] ), .B(\register_r[17][31] ), .C(
        \register_r[18][31] ), .D(\register_r[19][31] ), .S0(n2561), .S1(n2542), .Y(n2362) );
  MXI4X1 U1000 ( .A(\register_r[16][30] ), .B(\register_r[17][30] ), .C(
        \register_r[18][30] ), .D(\register_r[19][30] ), .S0(n2560), .S1(n2542), .Y(n2354) );
  MXI4X1 U1001 ( .A(\register_r[16][29] ), .B(\register_r[17][29] ), .C(
        \register_r[18][29] ), .D(\register_r[19][29] ), .S0(n2560), .S1(n2542), .Y(n2346) );
  MXI4X1 U1002 ( .A(\register_r[16][27] ), .B(\register_r[17][27] ), .C(
        \register_r[18][27] ), .D(\register_r[19][27] ), .S0(n2559), .S1(n2541), .Y(n2330) );
  MXI4X1 U1003 ( .A(\register_r[16][26] ), .B(\register_r[17][26] ), .C(
        \register_r[18][26] ), .D(\register_r[19][26] ), .S0(n2558), .S1(n2541), .Y(n2322) );
  MXI4X1 U1004 ( .A(\register_r[16][25] ), .B(\register_r[17][25] ), .C(
        \register_r[18][25] ), .D(\register_r[19][25] ), .S0(n2558), .S1(n2541), .Y(n2314) );
  MXI4X1 U1005 ( .A(\register_r[16][23] ), .B(\register_r[17][23] ), .C(
        \register_r[18][23] ), .D(\register_r[19][23] ), .S0(n2557), .S1(n2540), .Y(n2298) );
  MXI4X1 U1006 ( .A(\register_r[16][22] ), .B(\register_r[17][22] ), .C(
        \register_r[18][22] ), .D(\register_r[19][22] ), .S0(n2557), .S1(n2540), .Y(n2290) );
  MXI4X1 U1007 ( .A(\register_r[16][21] ), .B(\register_r[17][21] ), .C(
        \register_r[18][21] ), .D(\register_r[19][21] ), .S0(n2556), .S1(n2539), .Y(n2282) );
  MXI4X1 U1008 ( .A(\register_r[16][19] ), .B(\register_r[17][19] ), .C(
        \register_r[18][19] ), .D(\register_r[19][19] ), .S0(n2555), .S1(n2539), .Y(n2266) );
  MXI4X1 U1009 ( .A(\register_r[16][18] ), .B(\register_r[17][18] ), .C(
        \register_r[18][18] ), .D(\register_r[19][18] ), .S0(n2555), .S1(n2538), .Y(n2258) );
  MXI4X1 U1010 ( .A(\register_r[16][17] ), .B(\register_r[17][17] ), .C(
        \register_r[18][17] ), .D(\register_r[19][17] ), .S0(n2554), .S1(n2538), .Y(n2250) );
  MXI4X1 U1011 ( .A(\register_r[16][0] ), .B(\register_r[17][0] ), .C(
        \register_r[18][0] ), .D(\register_r[19][0] ), .S0(n2561), .S1(n2543), 
        .Y(n108) );
  MXI4X1 U1012 ( .A(\register_r[28][31] ), .B(\register_r[29][31] ), .C(
        \register_r[30][31] ), .D(\register_r[31][31] ), .S0(n2561), .S1(n2542), .Y(n2359) );
  MXI4X1 U1013 ( .A(\register_r[28][30] ), .B(\register_r[29][30] ), .C(
        \register_r[30][30] ), .D(\register_r[31][30] ), .S0(n2560), .S1(n2542), .Y(n2351) );
  MXI4X1 U1014 ( .A(\register_r[28][29] ), .B(\register_r[29][29] ), .C(
        \register_r[30][29] ), .D(\register_r[31][29] ), .S0(n2560), .S1(n2542), .Y(n2343) );
  MXI4X1 U1015 ( .A(\register_r[28][27] ), .B(\register_r[29][27] ), .C(
        \register_r[30][27] ), .D(\register_r[31][27] ), .S0(n2559), .S1(n2541), .Y(n2327) );
  MXI4X1 U1016 ( .A(\register_r[28][26] ), .B(\register_r[29][26] ), .C(
        \register_r[30][26] ), .D(\register_r[31][26] ), .S0(n2558), .S1(n2541), .Y(n2319) );
  MXI4X1 U1017 ( .A(\register_r[28][25] ), .B(\register_r[29][25] ), .C(
        \register_r[30][25] ), .D(\register_r[31][25] ), .S0(n2558), .S1(n2540), .Y(n2311) );
  MXI4X1 U1018 ( .A(\register_r[28][23] ), .B(\register_r[29][23] ), .C(
        \register_r[30][23] ), .D(\register_r[31][23] ), .S0(n2557), .S1(n2540), .Y(n2295) );
  MXI4X1 U1019 ( .A(\register_r[28][22] ), .B(\register_r[29][22] ), .C(
        \register_r[30][22] ), .D(\register_r[31][22] ), .S0(n2556), .S1(n2539), .Y(n2287) );
  MXI4X1 U1020 ( .A(\register_r[28][21] ), .B(\register_r[29][21] ), .C(
        \register_r[30][21] ), .D(\register_r[31][21] ), .S0(n2556), .S1(n2539), .Y(n2279) );
  MXI4X1 U1021 ( .A(\register_r[28][19] ), .B(\register_r[29][19] ), .C(
        \register_r[30][19] ), .D(\register_r[31][19] ), .S0(n2555), .S1(n2538), .Y(n2263) );
  MXI4X1 U1022 ( .A(\register_r[28][18] ), .B(\register_r[29][18] ), .C(
        \register_r[30][18] ), .D(\register_r[31][18] ), .S0(n2554), .S1(n2538), .Y(n2255) );
  MXI4X1 U1023 ( .A(\register_r[28][17] ), .B(\register_r[29][17] ), .C(
        \register_r[30][17] ), .D(\register_r[31][17] ), .S0(n2554), .S1(n2538), .Y(n2247) );
  MXI4X1 U1024 ( .A(r_12[15]), .B(r_13[15]), .C(\register_r[14][15] ), .D(
        \register_r[15][15] ), .S0(n2568), .S1(n2547), .Y(n2235) );
  MXI4X1 U1025 ( .A(r_12[14]), .B(r_13[14]), .C(\register_r[14][14] ), .D(
        \register_r[15][14] ), .S0(n2568), .S1(n2546), .Y(n2227) );
  MXI4X1 U1026 ( .A(r_12[13]), .B(r_13[13]), .C(\register_r[14][13] ), .D(
        \register_r[15][13] ), .S0(n2567), .S1(n2546), .Y(n2219) );
  MXI4X1 U1027 ( .A(r_12[11]), .B(r_13[11]), .C(\register_r[14][11] ), .D(
        \register_r[15][11] ), .S0(n2566), .S1(n2545), .Y(n2203) );
  MXI4X1 U1028 ( .A(r_12[10]), .B(r_13[10]), .C(\register_r[14][10] ), .D(
        \register_r[15][10] ), .S0(n2566), .S1(n2545), .Y(n2195) );
  MXI4X1 U1029 ( .A(r_12[9]), .B(r_13[9]), .C(\register_r[14][9] ), .D(
        \register_r[15][9] ), .S0(n2565), .S1(n2545), .Y(n2187) );
  MXI4X1 U1030 ( .A(r_12[7]), .B(r_13[7]), .C(\register_r[14][7] ), .D(
        \register_r[15][7] ), .S0(n2564), .S1(n2544), .Y(n2171) );
  MXI4X1 U1031 ( .A(r_12[6]), .B(r_13[6]), .C(\register_r[14][6] ), .D(
        \register_r[15][6] ), .S0(n2564), .S1(n2544), .Y(n2163) );
  MXI4X1 U1032 ( .A(r_12[5]), .B(r_13[5]), .C(\register_r[14][5] ), .D(
        \register_r[15][5] ), .S0(n2564), .S1(n2551), .Y(n2155) );
  MXI4X1 U1033 ( .A(r_12[3]), .B(r_13[3]), .C(\register_r[14][3] ), .D(
        \register_r[15][3] ), .S0(n2563), .S1(n2543), .Y(n2139) );
  MXI4X1 U1034 ( .A(r_12[2]), .B(r_13[2]), .C(\register_r[14][2] ), .D(
        \register_r[15][2] ), .S0(n2562), .S1(n2543), .Y(n2131) );
  MXI4X1 U1035 ( .A(r_12[1]), .B(r_13[1]), .C(\register_r[14][1] ), .D(
        \register_r[15][1] ), .S0(n2562), .S1(n2543), .Y(n2123) );
  MXI4X1 U1036 ( .A(\register_r[28][0] ), .B(\register_r[29][0] ), .C(
        \register_r[30][0] ), .D(\register_r[31][0] ), .S0(n2561), .S1(n2543), 
        .Y(n99) );
  MXI4X1 U1037 ( .A(\register_r[24][31] ), .B(\register_r[25][31] ), .C(
        \register_r[26][31] ), .D(\register_r[27][31] ), .S0(n2561), .S1(n2542), .Y(n2360) );
  MXI4X1 U1038 ( .A(\register_r[24][30] ), .B(\register_r[25][30] ), .C(
        \register_r[26][30] ), .D(\register_r[27][30] ), .S0(n2560), .S1(n2542), .Y(n2352) );
  MXI4X1 U1039 ( .A(\register_r[24][29] ), .B(\register_r[25][29] ), .C(
        \register_r[26][29] ), .D(\register_r[27][29] ), .S0(n2560), .S1(n2542), .Y(n2344) );
  MXI4X1 U1040 ( .A(\register_r[24][27] ), .B(\register_r[25][27] ), .C(
        \register_r[26][27] ), .D(\register_r[27][27] ), .S0(n2559), .S1(n2541), .Y(n2328) );
  MXI4X1 U1041 ( .A(\register_r[24][26] ), .B(\register_r[25][26] ), .C(
        \register_r[26][26] ), .D(\register_r[27][26] ), .S0(n2558), .S1(n2541), .Y(n2320) );
  MXI4X1 U1042 ( .A(\register_r[24][25] ), .B(\register_r[25][25] ), .C(
        \register_r[26][25] ), .D(\register_r[27][25] ), .S0(n2558), .S1(n2540), .Y(n2312) );
  MXI4X1 U1043 ( .A(\register_r[24][23] ), .B(\register_r[25][23] ), .C(
        \register_r[26][23] ), .D(\register_r[27][23] ), .S0(n2557), .S1(n2540), .Y(n2296) );
  MXI4X1 U1044 ( .A(\register_r[24][22] ), .B(\register_r[25][22] ), .C(
        \register_r[26][22] ), .D(\register_r[27][22] ), .S0(n2556), .S1(n2539), .Y(n2288) );
  MXI4X1 U1045 ( .A(\register_r[24][21] ), .B(\register_r[25][21] ), .C(
        \register_r[26][21] ), .D(\register_r[27][21] ), .S0(n2556), .S1(n2539), .Y(n2280) );
  MXI4X1 U1046 ( .A(\register_r[24][19] ), .B(\register_r[25][19] ), .C(
        \register_r[26][19] ), .D(\register_r[27][19] ), .S0(n2555), .S1(n2539), .Y(n2264) );
  MXI4X1 U1047 ( .A(\register_r[24][18] ), .B(\register_r[25][18] ), .C(
        \register_r[26][18] ), .D(\register_r[27][18] ), .S0(n2555), .S1(n2538), .Y(n2256) );
  MXI4X1 U1048 ( .A(\register_r[24][17] ), .B(\register_r[25][17] ), .C(
        \register_r[26][17] ), .D(\register_r[27][17] ), .S0(n2554), .S1(n2538), .Y(n2248) );
  MXI4X1 U1049 ( .A(\register_r[8][15] ), .B(\register_r[9][15] ), .C(
        \register_r[10][15] ), .D(\register_r[11][15] ), .S0(n2568), .S1(n2547), .Y(n2236) );
  MXI4X1 U1050 ( .A(\register_r[8][14] ), .B(\register_r[9][14] ), .C(
        \register_r[10][14] ), .D(\register_r[11][14] ), .S0(n2568), .S1(n2546), .Y(n2228) );
  MXI4X1 U1051 ( .A(\register_r[8][13] ), .B(\register_r[9][13] ), .C(
        \register_r[10][13] ), .D(\register_r[11][13] ), .S0(n2567), .S1(n2546), .Y(n2220) );
  MXI4X1 U1052 ( .A(\register_r[8][11] ), .B(\register_r[9][11] ), .C(
        \register_r[10][11] ), .D(\register_r[11][11] ), .S0(n2566), .S1(n2545), .Y(n2204) );
  MXI4X1 U1053 ( .A(\register_r[8][10] ), .B(\register_r[9][10] ), .C(
        \register_r[10][10] ), .D(\register_r[11][10] ), .S0(n2566), .S1(n2545), .Y(n2196) );
  MXI4X1 U1054 ( .A(\register_r[8][9] ), .B(\register_r[9][9] ), .C(
        \register_r[10][9] ), .D(\register_r[11][9] ), .S0(n2566), .S1(n2545), 
        .Y(n2188) );
  MXI4X1 U1055 ( .A(\register_r[8][7] ), .B(\register_r[9][7] ), .C(
        \register_r[10][7] ), .D(\register_r[11][7] ), .S0(n2565), .S1(n2544), 
        .Y(n2172) );
  MXI4X1 U1056 ( .A(\register_r[8][6] ), .B(\register_r[9][6] ), .C(
        \register_r[10][6] ), .D(\register_r[11][6] ), .S0(n2564), .S1(n2544), 
        .Y(n2164) );
  MXI4X1 U1057 ( .A(\register_r[8][5] ), .B(\register_r[9][5] ), .C(
        \register_r[10][5] ), .D(\register_r[11][5] ), .S0(n2564), .S1(n2551), 
        .Y(n2156) );
  MXI4X1 U1058 ( .A(\register_r[8][3] ), .B(\register_r[9][3] ), .C(
        \register_r[10][3] ), .D(\register_r[11][3] ), .S0(n2563), .S1(n2538), 
        .Y(n2140) );
  MXI4X1 U1059 ( .A(\register_r[8][2] ), .B(\register_r[9][2] ), .C(
        \register_r[10][2] ), .D(\register_r[11][2] ), .S0(n2562), .S1(n2543), 
        .Y(n2132) );
  MXI4X1 U1060 ( .A(\register_r[8][1] ), .B(\register_r[9][1] ), .C(
        \register_r[10][1] ), .D(\register_r[11][1] ), .S0(n2562), .S1(n2543), 
        .Y(n2124) );
  MXI4X1 U1061 ( .A(\register_r[24][0] ), .B(\register_r[25][0] ), .C(
        \register_r[26][0] ), .D(\register_r[27][0] ), .S0(n2561), .S1(n2543), 
        .Y(n102) );
  NAND4X1 U1062 ( .A(n126), .B(n127), .C(n128), .D(n129), .Y(n125) );
  XNOR2X1 U1063 ( .A(WriteReg[4]), .B(N11), .Y(n127) );
  XOR2X1 U1064 ( .A(n3442), .B(n3056), .Y(n128) );
  XOR2X1 U1065 ( .A(n3443), .B(N9), .Y(n126) );
  NAND4X1 U1066 ( .A(n133), .B(n134), .C(n135), .D(n136), .Y(n132) );
  XNOR2X1 U1067 ( .A(WriteReg[4]), .B(N6), .Y(n135) );
  XOR2X1 U1068 ( .A(n3442), .B(N5), .Y(n134) );
  XOR2X1 U1069 ( .A(n3443), .B(N4), .Y(n133) );
  CLKINVX1 U1070 ( .A(WriteReg[2]), .Y(n3443) );
  CLKINVX1 U1071 ( .A(WriteReg[3]), .Y(n3442) );
  CLKINVX1 U1072 ( .A(RegWrite), .Y(n3440) );
  NOR3X1 U1073 ( .A(n130), .B(n3440), .C(n131), .Y(n129) );
  XOR2X1 U1074 ( .A(WriteReg[1]), .B(N8), .Y(n130) );
  XOR2X1 U1075 ( .A(WriteReg[0]), .B(N7), .Y(n131) );
  NOR3X1 U1076 ( .A(n137), .B(n3440), .C(n138), .Y(n136) );
  XOR2X1 U1077 ( .A(WriteReg[1]), .B(N3), .Y(n137) );
  XOR2X1 U1078 ( .A(WriteReg[0]), .B(N2), .Y(n138) );
  MXI2X1 U1079 ( .A(n1067), .B(n2894), .S0(n3098), .Y(n2897) );
  NOR2BX1 U1080 ( .AN(n3075), .B(\register_r[3][31] ), .Y(n2894) );
  MX4X1 U1081 ( .A(n2789), .B(n2787), .C(n2788), .D(n2786), .S0(n3056), .S1(
        n3063), .Y(n2610) );
  MXI4X1 U1082 ( .A(\register_r[8][18] ), .B(\register_r[9][18] ), .C(
        \register_r[10][18] ), .D(\register_r[11][18] ), .S0(n3084), .S1(n3065), .Y(n2787) );
  MXI4X1 U1083 ( .A(r_12[18]), .B(r_13[18]), .C(\register_r[14][18] ), .D(
        \register_r[15][18] ), .S0(n3084), .S1(n3065), .Y(n2786) );
  MXI4X1 U1084 ( .A(\register_r[4][18] ), .B(\register_r[5][18] ), .C(
        \register_r[6][18] ), .D(\register_r[7][18] ), .S0(n3084), .S1(n3065), 
        .Y(n2788) );
  MX4X1 U1085 ( .A(n2781), .B(n2779), .C(n2780), .D(n2778), .S0(n3056), .S1(
        n3063), .Y(n2608) );
  MXI4X1 U1086 ( .A(\register_r[8][17] ), .B(\register_r[9][17] ), .C(
        \register_r[10][17] ), .D(\register_r[11][17] ), .S0(n3083), .S1(n3065), .Y(n2779) );
  MXI4X1 U1087 ( .A(r_12[17]), .B(r_13[17]), .C(\register_r[14][17] ), .D(
        \register_r[15][17] ), .S0(n3083), .S1(n3065), .Y(n2778) );
  MXI4X1 U1088 ( .A(\register_r[4][17] ), .B(\register_r[5][17] ), .C(
        \register_r[6][17] ), .D(\register_r[7][17] ), .S0(n3083), .S1(n3065), 
        .Y(n2780) );
  MX4X1 U1089 ( .A(n2773), .B(n2771), .C(n2772), .D(n2770), .S0(n3056), .S1(
        n3063), .Y(n2606) );
  MXI4X1 U1090 ( .A(\register_r[8][16] ), .B(\register_r[9][16] ), .C(
        \register_r[10][16] ), .D(\register_r[11][16] ), .S0(n3083), .S1(n3065), .Y(n2771) );
  MXI4X1 U1091 ( .A(r_12[16]), .B(r_13[16]), .C(\register_r[14][16] ), .D(
        \register_r[15][16] ), .S0(n3083), .S1(n3065), .Y(n2770) );
  MXI4X1 U1092 ( .A(\register_r[4][16] ), .B(\register_r[5][16] ), .C(
        \register_r[6][16] ), .D(\register_r[7][16] ), .S0(n3083), .S1(n3065), 
        .Y(n2772) );
  MX4X1 U1093 ( .A(n2893), .B(n2891), .C(n2892), .D(n2890), .S0(n3060), .S1(
        n3064), .Y(n2636) );
  MXI4X1 U1094 ( .A(\register_r[8][31] ), .B(\register_r[9][31] ), .C(
        \register_r[10][31] ), .D(\register_r[11][31] ), .S0(n3086), .S1(n3069), .Y(n2891) );
  MXI4X1 U1095 ( .A(r_12[31]), .B(r_13[31]), .C(\register_r[14][31] ), .D(
        \register_r[15][31] ), .S0(n3090), .S1(n3069), .Y(n2890) );
  NAND2X1 U1096 ( .A(n2898), .B(n2897), .Y(n2893) );
  MX4X1 U1097 ( .A(n2885), .B(n2883), .C(n2884), .D(n2882), .S0(n3060), .S1(
        n3063), .Y(n2634) );
  MXI4X1 U1098 ( .A(\register_r[8][30] ), .B(\register_r[9][30] ), .C(
        \register_r[10][30] ), .D(\register_r[11][30] ), .S0(n3089), .S1(n3068), .Y(n2883) );
  MXI4X1 U1099 ( .A(r_12[30]), .B(r_13[30]), .C(\register_r[14][30] ), .D(
        \register_r[15][30] ), .S0(n3089), .S1(n3068), .Y(n2882) );
  MXI4X1 U1100 ( .A(\register_r[4][30] ), .B(\register_r[5][30] ), .C(
        \register_r[6][30] ), .D(\register_r[7][30] ), .S0(n3090), .S1(n3068), 
        .Y(n2884) );
  MX4X1 U1101 ( .A(n2877), .B(n2875), .C(n2876), .D(n2874), .S0(n3060), .S1(
        n3063), .Y(n2632) );
  MXI4X1 U1102 ( .A(\register_r[8][29] ), .B(\register_r[9][29] ), .C(
        \register_r[10][29] ), .D(\register_r[11][29] ), .S0(n3089), .S1(n3068), .Y(n2875) );
  MXI4X1 U1103 ( .A(r_12[29]), .B(r_13[29]), .C(\register_r[14][29] ), .D(
        \register_r[15][29] ), .S0(n3089), .S1(n3068), .Y(n2874) );
  MXI4X1 U1104 ( .A(\register_r[4][29] ), .B(\register_r[5][29] ), .C(
        \register_r[6][29] ), .D(\register_r[7][29] ), .S0(n3089), .S1(n3068), 
        .Y(n2876) );
  MX4X1 U1105 ( .A(n2342), .B(n2340), .C(n2341), .D(n2339), .S0(n2533), .S1(
        n2537), .Y(n82) );
  MXI4X1 U1106 ( .A(\register_r[8][28] ), .B(\register_r[9][28] ), .C(
        \register_r[10][28] ), .D(\register_r[11][28] ), .S0(n2560), .S1(n2542), .Y(n2340) );
  MXI4X1 U1107 ( .A(r_12[28]), .B(r_13[28]), .C(\register_r[14][28] ), .D(
        \register_r[15][28] ), .S0(n2559), .S1(n2542), .Y(n2339) );
  MXI4X1 U1108 ( .A(\register_r[4][28] ), .B(\register_r[5][28] ), .C(
        \register_r[6][28] ), .D(\register_r[7][28] ), .S0(n2560), .S1(n2542), 
        .Y(n2341) );
  MX4X1 U1109 ( .A(n2869), .B(n2867), .C(n2868), .D(n2866), .S0(n3060), .S1(
        n3064), .Y(n2630) );
  MXI4X1 U1110 ( .A(\register_r[8][28] ), .B(\register_r[9][28] ), .C(
        \register_r[10][28] ), .D(\register_r[11][28] ), .S0(n3089), .S1(n3068), .Y(n2867) );
  MXI4X1 U1111 ( .A(r_12[28]), .B(r_13[28]), .C(\register_r[14][28] ), .D(
        \register_r[15][28] ), .S0(n3088), .S1(n3068), .Y(n2866) );
  MXI4X1 U1112 ( .A(\register_r[4][28] ), .B(\register_r[5][28] ), .C(
        \register_r[6][28] ), .D(\register_r[7][28] ), .S0(n3089), .S1(n3068), 
        .Y(n2868) );
  MX4X1 U1113 ( .A(n2829), .B(n2827), .C(n2828), .D(n2826), .S0(n3059), .S1(
        n3064), .Y(n2620) );
  MXI4X1 U1114 ( .A(\register_r[8][23] ), .B(\register_r[9][23] ), .C(
        \register_r[10][23] ), .D(\register_r[11][23] ), .S0(n3086), .S1(n3076), .Y(n2827) );
  MXI4X1 U1115 ( .A(r_12[23]), .B(r_13[23]), .C(\register_r[14][23] ), .D(
        \register_r[15][23] ), .S0(n3086), .S1(n3072), .Y(n2826) );
  MXI4X1 U1116 ( .A(\register_r[4][23] ), .B(\register_r[5][23] ), .C(
        \register_r[6][23] ), .D(\register_r[7][23] ), .S0(n3086), .S1(n3071), 
        .Y(n2828) );
  MX4X1 U1117 ( .A(n2821), .B(n2819), .C(n2820), .D(n2818), .S0(n3059), .S1(
        n3064), .Y(n2618) );
  MXI4X1 U1118 ( .A(\register_r[8][22] ), .B(\register_r[9][22] ), .C(
        \register_r[10][22] ), .D(\register_r[11][22] ), .S0(n3086), .S1(n3076), .Y(n2819) );
  MXI4X1 U1119 ( .A(r_12[22]), .B(r_13[22]), .C(\register_r[14][22] ), .D(
        \register_r[15][22] ), .S0(n3086), .S1(n3070), .Y(n2818) );
  MXI4X1 U1120 ( .A(\register_r[4][22] ), .B(\register_r[5][22] ), .C(
        \register_r[6][22] ), .D(\register_r[7][22] ), .S0(n3086), .S1(n3071), 
        .Y(n2820) );
  MX4X1 U1121 ( .A(n2813), .B(n2811), .C(n2812), .D(n2810), .S0(n3059), .S1(
        n3064), .Y(n2616) );
  MXI4X1 U1122 ( .A(\register_r[8][21] ), .B(\register_r[9][21] ), .C(
        \register_r[10][21] ), .D(\register_r[11][21] ), .S0(n3085), .S1(n3066), .Y(n2811) );
  MXI4X1 U1123 ( .A(r_12[21]), .B(r_13[21]), .C(\register_r[14][21] ), .D(
        \register_r[15][21] ), .S0(n3085), .S1(n3066), .Y(n2810) );
  MXI4X1 U1124 ( .A(\register_r[4][21] ), .B(\register_r[5][21] ), .C(
        \register_r[6][21] ), .D(\register_r[7][21] ), .S0(n3085), .S1(n3066), 
        .Y(n2812) );
  MX4X1 U1125 ( .A(n2805), .B(n2803), .C(n2804), .D(n2802), .S0(n3059), .S1(
        n3064), .Y(n2614) );
  MXI4X1 U1126 ( .A(\register_r[8][20] ), .B(\register_r[9][20] ), .C(
        \register_r[10][20] ), .D(\register_r[11][20] ), .S0(n3085), .S1(n3066), .Y(n2803) );
  MXI4X1 U1127 ( .A(r_12[20]), .B(r_13[20]), .C(\register_r[14][20] ), .D(
        \register_r[15][20] ), .S0(n3085), .S1(n3066), .Y(n2802) );
  MXI4X1 U1128 ( .A(\register_r[4][20] ), .B(\register_r[5][20] ), .C(
        \register_r[6][20] ), .D(\register_r[7][20] ), .S0(n3085), .S1(n3066), 
        .Y(n2804) );
  MX4X1 U1129 ( .A(n2853), .B(n2851), .C(n2852), .D(n2850), .S0(n3060), .S1(
        n3064), .Y(n2626) );
  MXI4X1 U1130 ( .A(\register_r[8][26] ), .B(\register_r[9][26] ), .C(
        \register_r[10][26] ), .D(\register_r[11][26] ), .S0(n3088), .S1(n3067), .Y(n2851) );
  MXI4X1 U1131 ( .A(r_12[26]), .B(r_13[26]), .C(\register_r[14][26] ), .D(
        \register_r[15][26] ), .S0(n3088), .S1(n3067), .Y(n2850) );
  MXI4X1 U1132 ( .A(\register_r[4][26] ), .B(\register_r[5][26] ), .C(
        \register_r[6][26] ), .D(\register_r[7][26] ), .S0(n3088), .S1(n3067), 
        .Y(n2852) );
  MX4X1 U1133 ( .A(n2861), .B(n2859), .C(n2860), .D(n2858), .S0(n3060), .S1(
        n3062), .Y(n2628) );
  MXI4X1 U1134 ( .A(\register_r[8][27] ), .B(\register_r[9][27] ), .C(
        \register_r[10][27] ), .D(\register_r[11][27] ), .S0(n3088), .S1(n3067), .Y(n2859) );
  MXI4X1 U1135 ( .A(r_12[27]), .B(r_13[27]), .C(\register_r[14][27] ), .D(
        \register_r[15][27] ), .S0(n3088), .S1(n3067), .Y(n2858) );
  MXI4X1 U1136 ( .A(\register_r[4][27] ), .B(\register_r[5][27] ), .C(
        \register_r[6][27] ), .D(\register_r[7][27] ), .S0(n3088), .S1(n3067), 
        .Y(n2860) );
  MX4X1 U1137 ( .A(n2845), .B(n2843), .C(n2844), .D(n2842), .S0(n3059), .S1(
        n3064), .Y(n2624) );
  MXI4X1 U1138 ( .A(\register_r[8][25] ), .B(\register_r[9][25] ), .C(
        \register_r[10][25] ), .D(\register_r[11][25] ), .S0(n3087), .S1(n3067), .Y(n2843) );
  MXI4X1 U1139 ( .A(r_12[25]), .B(r_13[25]), .C(\register_r[14][25] ), .D(
        \register_r[15][25] ), .S0(n3087), .S1(n3067), .Y(n2842) );
  MXI4X1 U1140 ( .A(\register_r[4][25] ), .B(\register_r[5][25] ), .C(
        \register_r[6][25] ), .D(\register_r[7][25] ), .S0(n3087), .S1(n3067), 
        .Y(n2844) );
  MX4X1 U1141 ( .A(n2837), .B(n2835), .C(n2836), .D(n2834), .S0(n3059), .S1(
        n3064), .Y(n2622) );
  MXI4X1 U1142 ( .A(\register_r[8][24] ), .B(\register_r[9][24] ), .C(
        \register_r[10][24] ), .D(\register_r[11][24] ), .S0(n3087), .S1(n3078), .Y(n2835) );
  MXI4X1 U1143 ( .A(r_12[24]), .B(r_13[24]), .C(\register_r[14][24] ), .D(
        \register_r[15][24] ), .S0(n3087), .S1(n3077), .Y(n2834) );
  MXI4X1 U1144 ( .A(\register_r[4][24] ), .B(\register_r[5][24] ), .C(
        \register_r[6][24] ), .D(\register_r[7][24] ), .S0(n3087), .S1(n3076), 
        .Y(n2836) );
  MX4X1 U1145 ( .A(n2310), .B(n2308), .C(n2309), .D(n2307), .S0(n2532), .S1(
        n2536), .Y(n63) );
  MXI4X1 U1146 ( .A(\register_r[8][24] ), .B(\register_r[9][24] ), .C(
        \register_r[10][24] ), .D(\register_r[11][24] ), .S0(n2558), .S1(n2540), .Y(n2308) );
  MXI4X1 U1147 ( .A(r_12[24]), .B(r_13[24]), .C(\register_r[14][24] ), .D(
        \register_r[15][24] ), .S0(n2558), .S1(n2540), .Y(n2307) );
  MXI4X1 U1148 ( .A(\register_r[4][24] ), .B(\register_r[5][24] ), .C(
        \register_r[6][24] ), .D(\register_r[7][24] ), .S0(n2558), .S1(n2540), 
        .Y(n2309) );
  MX4X1 U1149 ( .A(n2278), .B(n2276), .C(n2277), .D(n2275), .S0(n2532), .S1(
        n2536), .Y(n42) );
  MXI4X1 U1150 ( .A(\register_r[8][20] ), .B(\register_r[9][20] ), .C(
        \register_r[10][20] ), .D(\register_r[11][20] ), .S0(n2556), .S1(n2539), .Y(n2276) );
  MXI4X1 U1151 ( .A(r_12[20]), .B(r_13[20]), .C(\register_r[14][20] ), .D(
        \register_r[15][20] ), .S0(n2556), .S1(n2539), .Y(n2275) );
  MXI4X1 U1152 ( .A(\register_r[4][20] ), .B(\register_r[5][20] ), .C(
        \register_r[6][20] ), .D(\register_r[7][20] ), .S0(n2556), .S1(n2539), 
        .Y(n2277) );
  MX4X1 U1153 ( .A(n2246), .B(n2244), .C(n2245), .D(n2243), .S0(n2531), .S1(
        n2535), .Y(n34) );
  MXI4X1 U1154 ( .A(\register_r[8][16] ), .B(\register_r[9][16] ), .C(
        \register_r[10][16] ), .D(\register_r[11][16] ), .S0(n2554), .S1(n2538), .Y(n2244) );
  MXI4X1 U1155 ( .A(r_12[16]), .B(r_13[16]), .C(\register_r[14][16] ), .D(
        \register_r[15][16] ), .S0(n2554), .S1(n2538), .Y(n2243) );
  MXI4X1 U1156 ( .A(\register_r[4][16] ), .B(\register_r[5][16] ), .C(
        \register_r[6][16] ), .D(\register_r[7][16] ), .S0(n2554), .S1(n2538), 
        .Y(n2245) );
  MX4X1 U1157 ( .A(n2645), .B(n2643), .C(n2644), .D(n2642), .S0(n3058), .S1(
        n3061), .Y(n2574) );
  MXI4X1 U1158 ( .A(\register_r[8][0] ), .B(\register_r[9][0] ), .C(
        \register_r[10][0] ), .D(\register_r[11][0] ), .S0(n3090), .S1(n3069), 
        .Y(n2643) );
  MXI4X1 U1159 ( .A(r_12[0]), .B(r_13[0]), .C(\register_r[14][0] ), .D(
        \register_r[15][0] ), .S0(n3090), .S1(n3069), .Y(n2642) );
  MXI4X1 U1160 ( .A(\register_r[4][0] ), .B(\register_r[5][0] ), .C(
        \register_r[6][0] ), .D(\register_r[7][0] ), .S0(n3090), .S1(n3069), 
        .Y(n2644) );
  MX4X1 U1161 ( .A(n2665), .B(n2663), .C(n2664), .D(n2662), .S0(n3057), .S1(
        n3062), .Y(n2581) );
  MXI4X1 U1162 ( .A(\register_r[16][3] ), .B(\register_r[17][3] ), .C(
        \register_r[18][3] ), .D(\register_r[19][3] ), .S0(n3081), .S1(n3070), 
        .Y(n2665) );
  MXI4X1 U1163 ( .A(\register_r[24][3] ), .B(\register_r[25][3] ), .C(
        \register_r[26][3] ), .D(\register_r[27][3] ), .S0(n3091), .S1(n3070), 
        .Y(n2663) );
  MXI4X1 U1164 ( .A(\register_r[28][3] ), .B(\register_r[29][3] ), .C(
        \register_r[30][3] ), .D(\register_r[31][3] ), .S0(n3091), .S1(n3070), 
        .Y(n2662) );
  MX4X1 U1165 ( .A(n2657), .B(n2655), .C(n2656), .D(n2654), .S0(n3057), .S1(
        n3062), .Y(n2579) );
  MXI4X1 U1166 ( .A(\register_r[16][2] ), .B(\register_r[17][2] ), .C(
        \register_r[18][2] ), .D(\register_r[19][2] ), .S0(n3091), .S1(n3069), 
        .Y(n2657) );
  MXI4X1 U1167 ( .A(\register_r[24][2] ), .B(\register_r[25][2] ), .C(
        \register_r[26][2] ), .D(\register_r[27][2] ), .S0(n3091), .S1(n3069), 
        .Y(n2655) );
  MXI4X1 U1168 ( .A(\register_r[28][2] ), .B(\register_r[29][2] ), .C(
        \register_r[30][2] ), .D(\register_r[31][2] ), .S0(n3091), .S1(n3069), 
        .Y(n2654) );
  MX4X1 U1169 ( .A(n2697), .B(n2695), .C(n2696), .D(n2694), .S0(n3057), .S1(
        n3062), .Y(n2589) );
  MXI4X1 U1170 ( .A(\register_r[16][7] ), .B(\register_r[17][7] ), .C(
        \register_r[18][7] ), .D(\register_r[19][7] ), .S0(n3092), .S1(n3071), 
        .Y(n2697) );
  MXI4X1 U1171 ( .A(\register_r[24][7] ), .B(\register_r[25][7] ), .C(
        \register_r[26][7] ), .D(\register_r[27][7] ), .S0(n3092), .S1(n3071), 
        .Y(n2695) );
  MXI4X1 U1172 ( .A(\register_r[28][7] ), .B(\register_r[29][7] ), .C(
        \register_r[30][7] ), .D(\register_r[31][7] ), .S0(n3092), .S1(n3071), 
        .Y(n2694) );
  MX4X1 U1173 ( .A(n2689), .B(n2687), .C(n2688), .D(n2686), .S0(n3057), .S1(
        n3062), .Y(n2587) );
  MXI4X1 U1174 ( .A(\register_r[16][6] ), .B(\register_r[17][6] ), .C(
        \register_r[18][6] ), .D(\register_r[19][6] ), .S0(n3092), .S1(n3071), 
        .Y(n2689) );
  MXI4X1 U1175 ( .A(\register_r[24][6] ), .B(\register_r[25][6] ), .C(
        \register_r[26][6] ), .D(\register_r[27][6] ), .S0(n3092), .S1(n3071), 
        .Y(n2687) );
  MXI4X1 U1176 ( .A(\register_r[28][6] ), .B(\register_r[29][6] ), .C(
        \register_r[30][6] ), .D(\register_r[31][6] ), .S0(n3092), .S1(n3070), 
        .Y(n2686) );
  MX4X1 U1177 ( .A(n2681), .B(n2679), .C(n2680), .D(n2678), .S0(n3057), .S1(
        n3062), .Y(n2585) );
  MXI4X1 U1178 ( .A(\register_r[16][5] ), .B(\register_r[17][5] ), .C(
        \register_r[18][5] ), .D(\register_r[19][5] ), .S0(n3081), .S1(n3070), 
        .Y(n2681) );
  MXI4X1 U1179 ( .A(\register_r[24][5] ), .B(\register_r[25][5] ), .C(
        \register_r[26][5] ), .D(\register_r[27][5] ), .S0(n3081), .S1(n3070), 
        .Y(n2679) );
  MXI4X1 U1180 ( .A(\register_r[28][5] ), .B(\register_r[29][5] ), .C(
        \register_r[30][5] ), .D(\register_r[31][5] ), .S0(n3081), .S1(n3070), 
        .Y(n2678) );
  MX4X1 U1181 ( .A(n2673), .B(n2671), .C(n2672), .D(n2670), .S0(n3057), .S1(
        n3062), .Y(n2583) );
  MXI4X1 U1182 ( .A(\register_r[16][4] ), .B(\register_r[17][4] ), .C(
        \register_r[18][4] ), .D(\register_r[19][4] ), .S0(n3092), .S1(n3070), 
        .Y(n2673) );
  MXI4X1 U1183 ( .A(\register_r[24][4] ), .B(\register_r[25][4] ), .C(
        \register_r[26][4] ), .D(\register_r[27][4] ), .S0(n3085), .S1(n3070), 
        .Y(n2671) );
  MXI4X1 U1184 ( .A(\register_r[28][4] ), .B(\register_r[29][4] ), .C(
        \register_r[30][4] ), .D(\register_r[31][4] ), .S0(n3081), .S1(n3070), 
        .Y(n2670) );
  MX4X1 U1185 ( .A(n2729), .B(n2727), .C(n2728), .D(n2726), .S0(n3058), .S1(
        n3061), .Y(n2597) );
  MXI4X1 U1186 ( .A(\register_r[16][11] ), .B(\register_r[17][11] ), .C(
        \register_r[18][11] ), .D(\register_r[19][11] ), .S0(n3094), .S1(n3072), .Y(n2729) );
  MXI4X1 U1187 ( .A(\register_r[24][11] ), .B(\register_r[25][11] ), .C(
        \register_r[26][11] ), .D(\register_r[27][11] ), .S0(n3094), .S1(n3072), .Y(n2727) );
  MXI4X1 U1188 ( .A(\register_r[28][11] ), .B(\register_r[29][11] ), .C(
        \register_r[30][11] ), .D(\register_r[31][11] ), .S0(n3094), .S1(n3072), .Y(n2726) );
  MX4X1 U1189 ( .A(n2721), .B(n2719), .C(n2720), .D(n2718), .S0(n3058), .S1(
        n3061), .Y(n2595) );
  MXI4X1 U1190 ( .A(\register_r[16][10] ), .B(\register_r[17][10] ), .C(
        \register_r[18][10] ), .D(\register_r[19][10] ), .S0(n3094), .S1(n3072), .Y(n2721) );
  MXI4X1 U1191 ( .A(\register_r[24][10] ), .B(\register_r[25][10] ), .C(
        \register_r[26][10] ), .D(\register_r[27][10] ), .S0(n3094), .S1(n3072), .Y(n2719) );
  MXI4X1 U1192 ( .A(\register_r[28][10] ), .B(\register_r[29][10] ), .C(
        \register_r[30][10] ), .D(\register_r[31][10] ), .S0(n3094), .S1(n3072), .Y(n2718) );
  MX4X1 U1193 ( .A(n2713), .B(n2711), .C(n2712), .D(n2710), .S0(n3058), .S1(
        n3061), .Y(n2593) );
  MXI4X1 U1194 ( .A(\register_r[16][9] ), .B(\register_r[17][9] ), .C(
        \register_r[18][9] ), .D(\register_r[19][9] ), .S0(n3093), .S1(n3072), 
        .Y(n2713) );
  MXI4X1 U1195 ( .A(\register_r[24][9] ), .B(\register_r[25][9] ), .C(
        \register_r[26][9] ), .D(\register_r[27][9] ), .S0(n3093), .S1(n3072), 
        .Y(n2711) );
  MXI4X1 U1196 ( .A(\register_r[28][9] ), .B(\register_r[29][9] ), .C(
        \register_r[30][9] ), .D(\register_r[31][9] ), .S0(n3093), .S1(n3071), 
        .Y(n2710) );
  MX4X1 U1197 ( .A(n2705), .B(n2703), .C(n2704), .D(n2702), .S0(n3058), .S1(
        n3064), .Y(n2591) );
  MXI4X1 U1198 ( .A(\register_r[16][8] ), .B(\register_r[17][8] ), .C(
        \register_r[18][8] ), .D(\register_r[19][8] ), .S0(n3093), .S1(n3071), 
        .Y(n2705) );
  MXI4X1 U1199 ( .A(\register_r[24][8] ), .B(\register_r[25][8] ), .C(
        \register_r[26][8] ), .D(\register_r[27][8] ), .S0(n3093), .S1(n3071), 
        .Y(n2703) );
  MXI4X1 U1200 ( .A(\register_r[28][8] ), .B(\register_r[29][8] ), .C(
        \register_r[30][8] ), .D(\register_r[31][8] ), .S0(n3096), .S1(n3074), 
        .Y(n2702) );
  MX4X1 U1201 ( .A(n2761), .B(n2759), .C(n2760), .D(n2758), .S0(n3056), .S1(
        n3063), .Y(n2605) );
  MXI4X1 U1202 ( .A(\register_r[16][15] ), .B(\register_r[17][15] ), .C(
        \register_r[18][15] ), .D(\register_r[19][15] ), .S0(n3096), .S1(n3073), .Y(n2761) );
  MXI4X1 U1203 ( .A(\register_r[24][15] ), .B(\register_r[25][15] ), .C(
        \register_r[26][15] ), .D(\register_r[27][15] ), .S0(n3096), .S1(n3073), .Y(n2759) );
  MXI4X1 U1204 ( .A(\register_r[28][15] ), .B(\register_r[29][15] ), .C(
        \register_r[30][15] ), .D(\register_r[31][15] ), .S0(n3096), .S1(n3073), .Y(n2758) );
  MX4X1 U1205 ( .A(n2753), .B(n2751), .C(n2752), .D(n2750), .S0(n3056), .S1(
        n3063), .Y(n2603) );
  MXI4X1 U1206 ( .A(\register_r[16][14] ), .B(\register_r[17][14] ), .C(
        \register_r[18][14] ), .D(\register_r[19][14] ), .S0(n3096), .S1(n3073), .Y(n2753) );
  MXI4X1 U1207 ( .A(\register_r[24][14] ), .B(\register_r[25][14] ), .C(
        \register_r[26][14] ), .D(\register_r[27][14] ), .S0(n3096), .S1(n3073), .Y(n2751) );
  MXI4X1 U1208 ( .A(\register_r[28][14] ), .B(\register_r[29][14] ), .C(
        \register_r[30][14] ), .D(\register_r[31][14] ), .S0(n3095), .S1(n3073), .Y(n2750) );
  MX4X1 U1209 ( .A(n2745), .B(n2743), .C(n2744), .D(n2742), .S0(n3058), .S1(
        n3061), .Y(n2601) );
  MXI4X1 U1210 ( .A(\register_r[16][13] ), .B(\register_r[17][13] ), .C(
        \register_r[18][13] ), .D(\register_r[19][13] ), .S0(n3095), .S1(n3073), .Y(n2745) );
  MXI4X1 U1211 ( .A(\register_r[24][13] ), .B(\register_r[25][13] ), .C(
        \register_r[26][13] ), .D(\register_r[27][13] ), .S0(n3095), .S1(n3073), .Y(n2743) );
  MXI4X1 U1212 ( .A(\register_r[28][13] ), .B(\register_r[29][13] ), .C(
        \register_r[30][13] ), .D(\register_r[31][13] ), .S0(n3095), .S1(n3073), .Y(n2742) );
  MX4X1 U1213 ( .A(n2737), .B(n2735), .C(n2736), .D(n2734), .S0(n3058), .S1(
        n3061), .Y(n2599) );
  MXI4X1 U1214 ( .A(\register_r[16][12] ), .B(\register_r[17][12] ), .C(
        \register_r[18][12] ), .D(\register_r[19][12] ), .S0(n3095), .S1(n3073), .Y(n2737) );
  MXI4X1 U1215 ( .A(\register_r[24][12] ), .B(\register_r[25][12] ), .C(
        \register_r[26][12] ), .D(\register_r[27][12] ), .S0(n3095), .S1(n3072), .Y(n2735) );
  MXI4X1 U1216 ( .A(\register_r[28][12] ), .B(\register_r[29][12] ), .C(
        \register_r[30][12] ), .D(\register_r[31][12] ), .S0(n3095), .S1(n3072), .Y(n2734) );
  MX4X1 U1217 ( .A(n2210), .B(n2208), .C(n2209), .D(n2207), .S0(n2530), .S1(
        n2534), .Y(n27) );
  MXI4X1 U1218 ( .A(\register_r[16][12] ), .B(\register_r[17][12] ), .C(
        \register_r[18][12] ), .D(\register_r[19][12] ), .S0(n2567), .S1(n2546), .Y(n2210) );
  MXI4X1 U1219 ( .A(\register_r[24][12] ), .B(\register_r[25][12] ), .C(
        \register_r[26][12] ), .D(\register_r[27][12] ), .S0(n2567), .S1(n2545), .Y(n2208) );
  MXI4X1 U1220 ( .A(\register_r[28][12] ), .B(\register_r[29][12] ), .C(
        \register_r[30][12] ), .D(\register_r[31][12] ), .S0(n2567), .S1(n2545), .Y(n2207) );
  MX4X1 U1221 ( .A(n2178), .B(n2176), .C(n2177), .D(n2175), .S0(n2530), .S1(
        n2534), .Y(n19) );
  MXI4X1 U1222 ( .A(\register_r[16][8] ), .B(\register_r[17][8] ), .C(
        \register_r[18][8] ), .D(\register_r[19][8] ), .S0(n2565), .S1(n2544), 
        .Y(n2178) );
  MXI4X1 U1223 ( .A(\register_r[24][8] ), .B(\register_r[25][8] ), .C(
        \register_r[26][8] ), .D(\register_r[27][8] ), .S0(n2565), .S1(n2544), 
        .Y(n2176) );
  MXI4X1 U1224 ( .A(\register_r[28][8] ), .B(\register_r[29][8] ), .C(
        \register_r[30][8] ), .D(\register_r[31][8] ), .S0(n2568), .S1(n2547), 
        .Y(n2175) );
  MX4X1 U1225 ( .A(n2146), .B(n2144), .C(n2145), .D(n2143), .S0(n2529), .S1(
        n2535), .Y(n11) );
  MXI4X1 U1226 ( .A(\register_r[16][4] ), .B(\register_r[17][4] ), .C(
        \register_r[18][4] ), .D(\register_r[19][4] ), .S0(n2563), .S1(n2544), 
        .Y(n2146) );
  MXI4X1 U1227 ( .A(\register_r[24][4] ), .B(\register_r[25][4] ), .C(
        \register_r[26][4] ), .D(\register_r[27][4] ), .S0(n2563), .S1(n2548), 
        .Y(n2144) );
  MXI4X1 U1228 ( .A(\register_r[28][4] ), .B(\register_r[29][4] ), .C(
        \register_r[30][4] ), .D(\register_r[31][4] ), .S0(n2563), .S1(n2551), 
        .Y(n2143) );
  MX4X1 U1229 ( .A(n2649), .B(n2647), .C(n2648), .D(n2646), .S0(n3059), .S1(
        n3061), .Y(n2577) );
  MXI4X1 U1230 ( .A(\register_r[24][1] ), .B(\register_r[25][1] ), .C(
        \register_r[26][1] ), .D(\register_r[27][1] ), .S0(n3090), .S1(n3069), 
        .Y(n2647) );
  MXI4X1 U1231 ( .A(\register_r[16][1] ), .B(\register_r[17][1] ), .C(
        \register_r[18][1] ), .D(\register_r[19][1] ), .S0(n3091), .S1(n3069), 
        .Y(n2649) );
  MXI4X1 U1232 ( .A(\register_r[28][1] ), .B(\register_r[29][1] ), .C(
        \register_r[30][1] ), .D(\register_r[31][1] ), .S0(n3090), .S1(n3069), 
        .Y(n2646) );
  NOR2BX1 U1233 ( .AN(n3074), .B(\register_r[3][18] ), .Y(n2959) );
  NOR2BX1 U1234 ( .AN(n3074), .B(\register_r[3][17] ), .Y(n2964) );
  NOR2BX1 U1235 ( .AN(n3074), .B(\register_r[3][16] ), .Y(n2969) );
  NOR2BX1 U1236 ( .AN(n3075), .B(\register_r[3][30] ), .Y(n2899) );
  NOR2BX1 U1237 ( .AN(n3075), .B(\register_r[3][29] ), .Y(n2904) );
  NOR2BX1 U1238 ( .AN(n2548), .B(\register_r[3][28] ), .Y(n2382) );
  NOR2BX1 U1239 ( .AN(n3075), .B(\register_r[3][28] ), .Y(n2909) );
  NOR2BX1 U1240 ( .AN(n3074), .B(\register_r[3][23] ), .Y(n2934) );
  NOR2BX1 U1241 ( .AN(n3074), .B(\register_r[3][22] ), .Y(n2939) );
  NOR2BX1 U1242 ( .AN(n3074), .B(\register_r[3][21] ), .Y(n2944) );
  NOR2BX1 U1243 ( .AN(n3074), .B(\register_r[3][20] ), .Y(n2949) );
  NOR2BX1 U1244 ( .AN(n3075), .B(\register_r[3][26] ), .Y(n2919) );
  NOR2BX1 U1245 ( .AN(n3075), .B(\register_r[3][27] ), .Y(n2914) );
  NOR2BX1 U1246 ( .AN(n3075), .B(\register_r[3][25] ), .Y(n2924) );
  NOR2BX1 U1247 ( .AN(n3074), .B(\register_r[3][24] ), .Y(n2929) );
  NOR2BX1 U1248 ( .AN(n3075), .B(\register_r[3][3] ), .Y(n3034) );
  NOR2BX1 U1249 ( .AN(n3075), .B(\register_r[3][2] ), .Y(n3039) );
  NOR2BX1 U1250 ( .AN(n3075), .B(\register_r[3][1] ), .Y(n3044) );
  NOR2BX1 U1251 ( .AN(n3075), .B(\register_r[3][0] ), .Y(n3049) );
  NOR2BX1 U1252 ( .AN(n3074), .B(\register_r[3][7] ), .Y(n3014) );
  NOR2BX1 U1253 ( .AN(n3075), .B(\register_r[3][6] ), .Y(n3019) );
  NOR2BX1 U1254 ( .AN(n3074), .B(\register_r[3][5] ), .Y(n3024) );
  NOR2BX1 U1255 ( .AN(n3075), .B(\register_r[3][4] ), .Y(n3029) );
  NOR2BX1 U1256 ( .AN(n3074), .B(\register_r[3][11] ), .Y(n2994) );
  NOR2BX1 U1257 ( .AN(n3074), .B(\register_r[3][10] ), .Y(n2999) );
  NOR2BX1 U1258 ( .AN(n3074), .B(\register_r[3][9] ), .Y(n3004) );
  NOR2BX1 U1259 ( .AN(n3074), .B(\register_r[3][8] ), .Y(n3009) );
  NOR2BX1 U1260 ( .AN(n3074), .B(\register_r[3][15] ), .Y(n2974) );
  NOR2BX1 U1261 ( .AN(n3074), .B(\register_r[3][14] ), .Y(n2979) );
  NOR2BX1 U1262 ( .AN(n3074), .B(\register_r[3][13] ), .Y(n2984) );
  NOR2BX1 U1263 ( .AN(n3075), .B(\register_r[3][12] ), .Y(n2989) );
  NOR2BX1 U1264 ( .AN(n2547), .B(\register_r[3][24] ), .Y(n2402) );
  NOR2BX1 U1265 ( .AN(n2547), .B(\register_r[3][20] ), .Y(n2422) );
  NOR2BX1 U1266 ( .AN(n2547), .B(\register_r[3][16] ), .Y(n2442) );
  NOR2BX1 U1267 ( .AN(n2548), .B(\register_r[3][12] ), .Y(n2462) );
  NOR2BX1 U1268 ( .AN(n2547), .B(\register_r[3][8] ), .Y(n2482) );
  NOR2BX1 U1269 ( .AN(n2548), .B(\register_r[3][4] ), .Y(n2502) );
  NOR2X1 U1270 ( .A(n2369), .B(n2368), .Y(n2371) );
  NOR2X1 U1271 ( .A(n2542), .B(\register_r[1][31] ), .Y(n2369) );
  NOR2X1 U1272 ( .A(n2549), .B(n2573), .Y(n2368) );
  NOR2X1 U1273 ( .A(n2896), .B(n2895), .Y(n2898) );
  NOR2X1 U1274 ( .A(n3078), .B(\register_r[1][31] ), .Y(n2896) );
  NOR2X1 U1275 ( .A(n3078), .B(n3101), .Y(n2895) );
  NOR2X1 U1276 ( .A(n3077), .B(\register_r[1][26] ), .Y(n2921) );
  NOR2X1 U1277 ( .A(n2549), .B(\register_r[1][26] ), .Y(n2394) );
  NAND2X1 U1278 ( .A(n3048), .B(n3047), .Y(n2653) );
  NOR2X1 U1279 ( .A(n3046), .B(n3045), .Y(n3048) );
  MXI2X1 U1280 ( .A(n1097), .B(n3044), .S0(n3096), .Y(n3047) );
  NOR2X1 U1281 ( .A(n3071), .B(\register_r[1][1] ), .Y(n3046) );
  NAND2X1 U1282 ( .A(n2963), .B(n2962), .Y(n2789) );
  NOR2X1 U1283 ( .A(n2961), .B(n2960), .Y(n2963) );
  MXI2X1 U1284 ( .A(n1080), .B(n2959), .S0(n3098), .Y(n2962) );
  NOR2X1 U1285 ( .A(n3079), .B(\register_r[1][18] ), .Y(n2961) );
  NAND2X1 U1286 ( .A(n2968), .B(n2967), .Y(n2781) );
  NOR2X1 U1287 ( .A(n2966), .B(n2965), .Y(n2968) );
  MXI2X1 U1288 ( .A(n1081), .B(n2964), .S0(n3098), .Y(n2967) );
  NOR2X1 U1289 ( .A(n3076), .B(\register_r[1][17] ), .Y(n2966) );
  NAND2X1 U1290 ( .A(n2973), .B(n2972), .Y(n2773) );
  NOR2X1 U1291 ( .A(n2971), .B(n2970), .Y(n2973) );
  MXI2X1 U1292 ( .A(n1082), .B(n2969), .S0(n3098), .Y(n2972) );
  NOR2X1 U1293 ( .A(n3073), .B(\register_r[1][16] ), .Y(n2971) );
  NAND2X1 U1294 ( .A(n2908), .B(n2907), .Y(n2877) );
  NOR2X1 U1295 ( .A(n2906), .B(n2905), .Y(n2908) );
  MXI2X1 U1296 ( .A(n1069), .B(n2904), .S0(n3098), .Y(n2907) );
  NOR2X1 U1297 ( .A(n3078), .B(\register_r[1][29] ), .Y(n2906) );
  NAND2X1 U1298 ( .A(n2938), .B(n2937), .Y(n2829) );
  NOR2X1 U1299 ( .A(n2936), .B(n2935), .Y(n2938) );
  MXI2X1 U1300 ( .A(n1075), .B(n2934), .S0(n3098), .Y(n2937) );
  NOR2X1 U1301 ( .A(n3077), .B(\register_r[1][23] ), .Y(n2936) );
  NAND2X1 U1302 ( .A(n2943), .B(n2942), .Y(n2821) );
  NOR2X1 U1303 ( .A(n2941), .B(n2940), .Y(n2943) );
  MXI2X1 U1304 ( .A(n1076), .B(n2939), .S0(n3098), .Y(n2942) );
  NOR2X1 U1305 ( .A(n3077), .B(\register_r[1][22] ), .Y(n2941) );
  NAND2X1 U1306 ( .A(n2948), .B(n2947), .Y(n2813) );
  NOR2X1 U1307 ( .A(n2946), .B(n2945), .Y(n2948) );
  MXI2X1 U1308 ( .A(n1077), .B(n2944), .S0(n3098), .Y(n2947) );
  NOR2X1 U1309 ( .A(n3077), .B(\register_r[1][21] ), .Y(n2946) );
  NAND2X1 U1310 ( .A(n2953), .B(n2952), .Y(n2805) );
  NOR2X1 U1311 ( .A(n2951), .B(n2950), .Y(n2953) );
  MXI2X1 U1312 ( .A(n1078), .B(n2949), .S0(n3098), .Y(n2952) );
  NOR2X1 U1313 ( .A(n3077), .B(\register_r[1][20] ), .Y(n2951) );
  NAND2X1 U1314 ( .A(n2923), .B(n2922), .Y(n2853) );
  NOR2X1 U1315 ( .A(n2921), .B(n2920), .Y(n2923) );
  MXI2X1 U1316 ( .A(n1072), .B(n2919), .S0(n3098), .Y(n2922) );
  NOR2X1 U1317 ( .A(n3078), .B(n3100), .Y(n2920) );
  NAND2X1 U1318 ( .A(n2933), .B(n2932), .Y(n2837) );
  NOR2X1 U1319 ( .A(n2931), .B(n2930), .Y(n2933) );
  MXI2X1 U1320 ( .A(n1074), .B(n2929), .S0(n3098), .Y(n2932) );
  NOR2X1 U1321 ( .A(n3077), .B(\register_r[1][24] ), .Y(n2931) );
  NAND2X1 U1322 ( .A(n3038), .B(n3037), .Y(n2669) );
  NOR2X1 U1323 ( .A(n3036), .B(n3035), .Y(n3038) );
  MXI2X1 U1324 ( .A(n1095), .B(n3034), .S0(n3097), .Y(n3037) );
  NOR2X1 U1325 ( .A(n3076), .B(\register_r[1][3] ), .Y(n3036) );
  NAND2X1 U1326 ( .A(n3043), .B(n3042), .Y(n2661) );
  NOR2X1 U1327 ( .A(n3041), .B(n3040), .Y(n3043) );
  MXI2X1 U1328 ( .A(n1096), .B(n3039), .S0(n3097), .Y(n3042) );
  NOR2X1 U1329 ( .A(n3078), .B(\register_r[1][2] ), .Y(n3041) );
  NAND2X1 U1330 ( .A(n3018), .B(n3017), .Y(n2701) );
  NOR2X1 U1331 ( .A(n3016), .B(n3015), .Y(n3018) );
  MXI2X1 U1332 ( .A(n1091), .B(n3014), .S0(n3097), .Y(n3017) );
  NOR2X1 U1333 ( .A(n3076), .B(\register_r[1][7] ), .Y(n3016) );
  NAND2X1 U1334 ( .A(n3023), .B(n3022), .Y(n2693) );
  NOR2X1 U1335 ( .A(n3021), .B(n3020), .Y(n3023) );
  MXI2X1 U1336 ( .A(n1092), .B(n3019), .S0(n3097), .Y(n3022) );
  NOR2X1 U1337 ( .A(n3075), .B(\register_r[1][6] ), .Y(n3021) );
  NAND2X1 U1338 ( .A(n3028), .B(n3027), .Y(n2685) );
  NOR2X1 U1339 ( .A(n3026), .B(n3025), .Y(n3028) );
  MXI2X1 U1340 ( .A(n1093), .B(n3024), .S0(n3097), .Y(n3027) );
  NOR2X1 U1341 ( .A(n3076), .B(\register_r[1][5] ), .Y(n3026) );
  NAND2X1 U1342 ( .A(n3033), .B(n3032), .Y(n2677) );
  NOR2X1 U1343 ( .A(n3031), .B(n3030), .Y(n3033) );
  MXI2X1 U1344 ( .A(n1094), .B(n3029), .S0(n3097), .Y(n3032) );
  NOR2X1 U1345 ( .A(n3075), .B(\register_r[1][4] ), .Y(n3031) );
  NAND2X1 U1346 ( .A(n2998), .B(n2997), .Y(n2733) );
  NOR2X1 U1347 ( .A(n2996), .B(n2995), .Y(n2998) );
  MXI2X1 U1348 ( .A(n1087), .B(n2994), .S0(n3097), .Y(n2997) );
  NOR2X1 U1349 ( .A(n3078), .B(\register_r[1][11] ), .Y(n2996) );
  NAND2X1 U1350 ( .A(n3003), .B(n3002), .Y(n2725) );
  NOR2X1 U1351 ( .A(n3001), .B(n3000), .Y(n3003) );
  MXI2X1 U1352 ( .A(n1088), .B(n2999), .S0(n3097), .Y(n3002) );
  NOR2X1 U1353 ( .A(n3076), .B(\register_r[1][10] ), .Y(n3001) );
  NAND2X1 U1354 ( .A(n3008), .B(n3007), .Y(n2717) );
  NOR2X1 U1355 ( .A(n3006), .B(n3005), .Y(n3008) );
  MXI2X1 U1356 ( .A(n1089), .B(n3004), .S0(n3097), .Y(n3007) );
  NOR2X1 U1357 ( .A(n3076), .B(\register_r[1][9] ), .Y(n3006) );
  NAND2X1 U1358 ( .A(n3013), .B(n3012), .Y(n2709) );
  NOR2X1 U1359 ( .A(n3011), .B(n3010), .Y(n3013) );
  MXI2X1 U1360 ( .A(n1090), .B(n3009), .S0(n3097), .Y(n3012) );
  NOR2X1 U1361 ( .A(n3072), .B(\register_r[1][8] ), .Y(n3011) );
  NAND2X1 U1362 ( .A(n2978), .B(n2977), .Y(n2765) );
  NOR2X1 U1363 ( .A(n2976), .B(n2975), .Y(n2978) );
  MXI2X1 U1364 ( .A(n1083), .B(n2974), .S0(n3098), .Y(n2977) );
  NOR2X1 U1365 ( .A(n3079), .B(\register_r[1][15] ), .Y(n2976) );
  NAND2X1 U1366 ( .A(n2983), .B(n2982), .Y(n2757) );
  NOR2X1 U1367 ( .A(n2981), .B(n2980), .Y(n2983) );
  MXI2X1 U1368 ( .A(n1084), .B(n2979), .S0(n3097), .Y(n2982) );
  NOR2X1 U1369 ( .A(n3076), .B(\register_r[1][14] ), .Y(n2981) );
  NAND2X1 U1370 ( .A(n2988), .B(n2987), .Y(n2749) );
  NOR2X1 U1371 ( .A(n2986), .B(n2985), .Y(n2988) );
  MXI2X1 U1372 ( .A(n1085), .B(n2984), .S0(n3097), .Y(n2987) );
  NOR2X1 U1373 ( .A(n3077), .B(\register_r[1][13] ), .Y(n2986) );
  NAND2X1 U1374 ( .A(n2993), .B(n2992), .Y(n2741) );
  NOR2X1 U1375 ( .A(n2991), .B(n2990), .Y(n2993) );
  MXI2X1 U1376 ( .A(n1086), .B(n2989), .S0(n3097), .Y(n2992) );
  NOR2X1 U1377 ( .A(n3070), .B(\register_r[1][12] ), .Y(n2991) );
  NAND2X1 U1378 ( .A(n2406), .B(n2405), .Y(n2310) );
  NOR2X1 U1379 ( .A(n2404), .B(n2403), .Y(n2406) );
  MXI2X1 U1380 ( .A(n1074), .B(n2402), .S0(n2570), .Y(n2405) );
  NOR2X1 U1381 ( .A(n2539), .B(\register_r[1][24] ), .Y(n2404) );
  NAND2X1 U1382 ( .A(n2426), .B(n2425), .Y(n2278) );
  NOR2X1 U1383 ( .A(n2424), .B(n2423), .Y(n2426) );
  MXI2X1 U1384 ( .A(n1078), .B(n2422), .S0(n2570), .Y(n2425) );
  NOR2X1 U1385 ( .A(n2545), .B(\register_r[1][20] ), .Y(n2424) );
  NAND2X1 U1386 ( .A(n2446), .B(n2445), .Y(n2246) );
  NOR2X1 U1387 ( .A(n2444), .B(n2443), .Y(n2446) );
  MXI2X1 U1388 ( .A(n1082), .B(n2442), .S0(n2570), .Y(n2445) );
  NOR2X1 U1389 ( .A(n2543), .B(\register_r[1][16] ), .Y(n2444) );
  NAND2X1 U1390 ( .A(n2466), .B(n2465), .Y(n2214) );
  NOR2X1 U1391 ( .A(n2464), .B(n2463), .Y(n2466) );
  MXI2X1 U1392 ( .A(n1086), .B(n2462), .S0(n2569), .Y(n2465) );
  NOR2X1 U1393 ( .A(n2550), .B(\register_r[1][12] ), .Y(n2464) );
  NAND2X1 U1394 ( .A(n2486), .B(n2485), .Y(n2182) );
  NOR2X1 U1395 ( .A(n2484), .B(n2483), .Y(n2486) );
  MXI2X1 U1396 ( .A(n1090), .B(n2482), .S0(n2569), .Y(n2485) );
  NOR2X1 U1397 ( .A(n2550), .B(\register_r[1][8] ), .Y(n2484) );
  NAND2X1 U1398 ( .A(n2506), .B(n2505), .Y(n2150) );
  NOR2X1 U1399 ( .A(n2504), .B(n2503), .Y(n2506) );
  MXI2X1 U1400 ( .A(n1094), .B(n2502), .S0(n2569), .Y(n2505) );
  NOR2X1 U1401 ( .A(n2548), .B(\register_r[1][4] ), .Y(n2504) );
  NAND2X1 U1402 ( .A(n2903), .B(n2902), .Y(n2885) );
  NOR2X1 U1403 ( .A(n2901), .B(n2900), .Y(n2903) );
  MXI2X1 U1404 ( .A(n1068), .B(n2899), .S0(n3099), .Y(n2902) );
  NOR2X1 U1405 ( .A(n3078), .B(\register_r[1][30] ), .Y(n2901) );
  NAND2X1 U1406 ( .A(n2386), .B(n2385), .Y(n2342) );
  NOR2X1 U1407 ( .A(n2384), .B(n2383), .Y(n2386) );
  MXI2X1 U1408 ( .A(n1070), .B(n2382), .S0(n2571), .Y(n2385) );
  NOR2X1 U1409 ( .A(n2539), .B(\register_r[1][28] ), .Y(n2384) );
  NAND2X1 U1410 ( .A(n2913), .B(n2912), .Y(n2869) );
  NOR2X1 U1411 ( .A(n2911), .B(n2910), .Y(n2913) );
  MXI2X1 U1412 ( .A(n1070), .B(n2909), .S0(n3099), .Y(n2912) );
  NOR2X1 U1413 ( .A(n3078), .B(\register_r[1][28] ), .Y(n2911) );
  NAND2X1 U1414 ( .A(n2918), .B(n2917), .Y(n2861) );
  NOR2X1 U1415 ( .A(n2916), .B(n2915), .Y(n2918) );
  MXI2X1 U1416 ( .A(n1071), .B(n2914), .S0(n3099), .Y(n2917) );
  NOR2X1 U1417 ( .A(n3078), .B(\register_r[1][27] ), .Y(n2916) );
  NAND2X1 U1418 ( .A(n2928), .B(n2927), .Y(n2845) );
  NOR2X1 U1419 ( .A(n2926), .B(n2925), .Y(n2928) );
  MXI2X1 U1420 ( .A(n1073), .B(n2924), .S0(n3099), .Y(n2927) );
  NOR2X1 U1421 ( .A(n3077), .B(\register_r[1][25] ), .Y(n2926) );
  NAND2X1 U1422 ( .A(n3053), .B(n3052), .Y(n2645) );
  NOR2X1 U1423 ( .A(n3051), .B(n3050), .Y(n3053) );
  MXI2X1 U1424 ( .A(n1098), .B(n3049), .S0(n3099), .Y(n3052) );
  NOR2X1 U1425 ( .A(n3078), .B(\register_r[1][0] ), .Y(n3051) );
  MXI4X1 U1426 ( .A(\register_r[20][19] ), .B(\register_r[21][19] ), .C(
        \register_r[22][19] ), .D(\register_r[23][19] ), .S0(n3084), .S1(n3066), .Y(n2792) );
  MXI4X1 U1427 ( .A(\register_r[20][18] ), .B(\register_r[21][18] ), .C(
        \register_r[22][18] ), .D(\register_r[23][18] ), .S0(n3084), .S1(n3065), .Y(n2784) );
  MXI4X1 U1428 ( .A(\register_r[20][17] ), .B(\register_r[21][17] ), .C(
        \register_r[22][17] ), .D(\register_r[23][17] ), .S0(n3083), .S1(n3065), .Y(n2776) );
  MXI4X1 U1429 ( .A(\register_r[20][16] ), .B(\register_r[21][16] ), .C(
        \register_r[22][16] ), .D(\register_r[23][16] ), .S0(n3083), .S1(n3065), .Y(n2768) );
  MXI4X1 U1430 ( .A(\register_r[4][31] ), .B(\register_r[5][31] ), .C(
        \register_r[6][31] ), .D(\register_r[7][31] ), .S0(n3096), .S1(n3074), 
        .Y(n2892) );
  MXI4X1 U1431 ( .A(\register_r[20][31] ), .B(\register_r[21][31] ), .C(
        \register_r[22][31] ), .D(\register_r[23][31] ), .S0(n3090), .S1(n3068), .Y(n2888) );
  MXI4X1 U1432 ( .A(\register_r[20][30] ), .B(\register_r[21][30] ), .C(
        \register_r[22][30] ), .D(\register_r[23][30] ), .S0(n3089), .S1(n3068), .Y(n2880) );
  MXI4X1 U1433 ( .A(\register_r[20][29] ), .B(\register_r[21][29] ), .C(
        \register_r[22][29] ), .D(\register_r[23][29] ), .S0(n3089), .S1(n3068), .Y(n2872) );
  MXI4X1 U1434 ( .A(\register_r[20][28] ), .B(\register_r[21][28] ), .C(
        \register_r[22][28] ), .D(\register_r[23][28] ), .S0(n2559), .S1(n2541), .Y(n2337) );
  MXI4X1 U1435 ( .A(\register_r[20][28] ), .B(\register_r[21][28] ), .C(
        \register_r[22][28] ), .D(\register_r[23][28] ), .S0(n3088), .S1(n3067), .Y(n2864) );
  MXI4X1 U1436 ( .A(\register_r[20][23] ), .B(\register_r[21][23] ), .C(
        \register_r[22][23] ), .D(\register_r[23][23] ), .S0(n3086), .S1(n3071), .Y(n2824) );
  MXI4X1 U1437 ( .A(\register_r[20][22] ), .B(\register_r[21][22] ), .C(
        \register_r[22][22] ), .D(\register_r[23][22] ), .S0(n3085), .S1(n3070), .Y(n2816) );
  MXI4X1 U1438 ( .A(\register_r[20][21] ), .B(\register_r[21][21] ), .C(
        \register_r[22][21] ), .D(\register_r[23][21] ), .S0(n3085), .S1(n3066), .Y(n2808) );
  MXI4X1 U1439 ( .A(\register_r[20][20] ), .B(\register_r[21][20] ), .C(
        \register_r[22][20] ), .D(\register_r[23][20] ), .S0(n3085), .S1(n3066), .Y(n2800) );
  MXI4X1 U1440 ( .A(\register_r[20][26] ), .B(\register_r[21][26] ), .C(
        \register_r[22][26] ), .D(\register_r[23][26] ), .S0(n3087), .S1(n3067), .Y(n2848) );
  MXI4X1 U1441 ( .A(\register_r[20][27] ), .B(\register_r[21][27] ), .C(
        \register_r[22][27] ), .D(\register_r[23][27] ), .S0(n3088), .S1(n3067), .Y(n2856) );
  MXI4X1 U1442 ( .A(\register_r[20][25] ), .B(\register_r[21][25] ), .C(
        \register_r[22][25] ), .D(\register_r[23][25] ), .S0(n3087), .S1(n3067), .Y(n2840) );
  MXI4X1 U1443 ( .A(\register_r[20][24] ), .B(\register_r[21][24] ), .C(
        \register_r[22][24] ), .D(\register_r[23][24] ), .S0(n3086), .S1(n3076), .Y(n2832) );
  MXI4X1 U1444 ( .A(\register_r[20][3] ), .B(\register_r[21][3] ), .C(
        \register_r[22][3] ), .D(\register_r[23][3] ), .S0(n3091), .S1(n3070), 
        .Y(n2664) );
  MXI4X1 U1445 ( .A(\register_r[4][3] ), .B(\register_r[5][3] ), .C(
        \register_r[6][3] ), .D(\register_r[7][3] ), .S0(n3081), .S1(n3070), 
        .Y(n2668) );
  MXI4X1 U1446 ( .A(\register_r[20][2] ), .B(\register_r[21][2] ), .C(
        \register_r[22][2] ), .D(\register_r[23][2] ), .S0(n3091), .S1(n3069), 
        .Y(n2656) );
  MXI4X1 U1447 ( .A(\register_r[4][2] ), .B(\register_r[5][2] ), .C(
        \register_r[6][2] ), .D(\register_r[7][2] ), .S0(n3091), .S1(n3069), 
        .Y(n2660) );
  MXI4X1 U1448 ( .A(\register_r[20][1] ), .B(\register_r[21][1] ), .C(
        \register_r[22][1] ), .D(\register_r[23][1] ), .S0(n3091), .S1(n3069), 
        .Y(n2648) );
  MXI4X1 U1449 ( .A(\register_r[4][1] ), .B(\register_r[5][1] ), .C(
        \register_r[6][1] ), .D(\register_r[7][1] ), .S0(n3091), .S1(n3069), 
        .Y(n2652) );
  MXI4X1 U1450 ( .A(\register_r[20][0] ), .B(\register_r[21][0] ), .C(
        \register_r[22][0] ), .D(\register_r[23][0] ), .S0(n3090), .S1(n3069), 
        .Y(n2640) );
  MXI4X1 U1451 ( .A(\register_r[20][7] ), .B(\register_r[21][7] ), .C(
        \register_r[22][7] ), .D(\register_r[23][7] ), .S0(n3092), .S1(n3071), 
        .Y(n2696) );
  MXI4X1 U1452 ( .A(\register_r[4][7] ), .B(\register_r[5][7] ), .C(
        \register_r[6][7] ), .D(\register_r[7][7] ), .S0(n3093), .S1(n3071), 
        .Y(n2700) );
  MXI4X1 U1453 ( .A(\register_r[20][6] ), .B(\register_r[21][6] ), .C(
        \register_r[22][6] ), .D(\register_r[23][6] ), .S0(n3092), .S1(n3071), 
        .Y(n2688) );
  MXI4X1 U1454 ( .A(\register_r[4][6] ), .B(\register_r[5][6] ), .C(
        \register_r[6][6] ), .D(\register_r[7][6] ), .S0(n3092), .S1(n3071), 
        .Y(n2692) );
  MXI4X1 U1455 ( .A(\register_r[20][5] ), .B(\register_r[21][5] ), .C(
        \register_r[22][5] ), .D(\register_r[23][5] ), .S0(n3081), .S1(n3070), 
        .Y(n2680) );
  MXI4X1 U1456 ( .A(\register_r[4][5] ), .B(\register_r[5][5] ), .C(
        \register_r[6][5] ), .D(\register_r[7][5] ), .S0(n3092), .S1(n3070), 
        .Y(n2684) );
  MXI4X1 U1457 ( .A(\register_r[20][4] ), .B(\register_r[21][4] ), .C(
        \register_r[22][4] ), .D(\register_r[23][4] ), .S0(n3091), .S1(n3070), 
        .Y(n2672) );
  MXI4X1 U1458 ( .A(\register_r[4][4] ), .B(\register_r[5][4] ), .C(
        \register_r[6][4] ), .D(\register_r[7][4] ), .S0(n3095), .S1(n3070), 
        .Y(n2676) );
  MXI4X1 U1459 ( .A(\register_r[20][11] ), .B(\register_r[21][11] ), .C(
        \register_r[22][11] ), .D(\register_r[23][11] ), .S0(n3094), .S1(n3072), .Y(n2728) );
  MXI4X1 U1460 ( .A(\register_r[4][11] ), .B(\register_r[5][11] ), .C(
        \register_r[6][11] ), .D(\register_r[7][11] ), .S0(n3095), .S1(n3072), 
        .Y(n2732) );
  MXI4X1 U1461 ( .A(\register_r[20][10] ), .B(\register_r[21][10] ), .C(
        \register_r[22][10] ), .D(\register_r[23][10] ), .S0(n3094), .S1(n3072), .Y(n2720) );
  MXI4X1 U1462 ( .A(\register_r[4][10] ), .B(\register_r[5][10] ), .C(
        \register_r[6][10] ), .D(\register_r[7][10] ), .S0(n3094), .S1(n3072), 
        .Y(n2724) );
  MXI4X1 U1463 ( .A(\register_r[20][9] ), .B(\register_r[21][9] ), .C(
        \register_r[22][9] ), .D(\register_r[23][9] ), .S0(n3093), .S1(n3072), 
        .Y(n2712) );
  MXI4X1 U1464 ( .A(\register_r[4][9] ), .B(\register_r[5][9] ), .C(
        \register_r[6][9] ), .D(\register_r[7][9] ), .S0(n3094), .S1(n3072), 
        .Y(n2716) );
  MXI4X1 U1465 ( .A(\register_r[20][8] ), .B(\register_r[21][8] ), .C(
        \register_r[22][8] ), .D(\register_r[23][8] ), .S0(n3093), .S1(n3071), 
        .Y(n2704) );
  MXI4X1 U1466 ( .A(\register_r[4][8] ), .B(\register_r[5][8] ), .C(
        \register_r[6][8] ), .D(\register_r[7][8] ), .S0(n3093), .S1(n3071), 
        .Y(n2708) );
  MXI4X1 U1467 ( .A(\register_r[20][15] ), .B(\register_r[21][15] ), .C(
        \register_r[22][15] ), .D(\register_r[23][15] ), .S0(n3096), .S1(n3073), .Y(n2760) );
  MXI4X1 U1468 ( .A(\register_r[4][15] ), .B(\register_r[5][15] ), .C(
        \register_r[6][15] ), .D(\register_r[7][15] ), .S0(n3093), .S1(n3071), 
        .Y(n2764) );
  MXI4X1 U1469 ( .A(\register_r[20][14] ), .B(\register_r[21][14] ), .C(
        \register_r[22][14] ), .D(\register_r[23][14] ), .S0(n3096), .S1(n3073), .Y(n2752) );
  MXI4X1 U1470 ( .A(\register_r[4][14] ), .B(\register_r[5][14] ), .C(
        \register_r[6][14] ), .D(\register_r[7][14] ), .S0(n3096), .S1(n3073), 
        .Y(n2756) );
  MXI4X1 U1471 ( .A(\register_r[20][13] ), .B(\register_r[21][13] ), .C(
        \register_r[22][13] ), .D(\register_r[23][13] ), .S0(n3095), .S1(n3073), .Y(n2744) );
  MXI4X1 U1472 ( .A(\register_r[4][13] ), .B(\register_r[5][13] ), .C(
        \register_r[6][13] ), .D(\register_r[7][13] ), .S0(n3095), .S1(n3073), 
        .Y(n2748) );
  MXI4X1 U1473 ( .A(\register_r[20][12] ), .B(\register_r[21][12] ), .C(
        \register_r[22][12] ), .D(\register_r[23][12] ), .S0(n3095), .S1(n3073), .Y(n2736) );
  MXI4X1 U1474 ( .A(\register_r[4][12] ), .B(\register_r[5][12] ), .C(
        \register_r[6][12] ), .D(\register_r[7][12] ), .S0(n3093), .S1(n3071), 
        .Y(n2740) );
  MXI4X1 U1475 ( .A(\register_r[20][24] ), .B(\register_r[21][24] ), .C(
        \register_r[22][24] ), .D(\register_r[23][24] ), .S0(n2557), .S1(n2540), .Y(n2305) );
  MXI4X1 U1476 ( .A(\register_r[20][20] ), .B(\register_r[21][20] ), .C(
        \register_r[22][20] ), .D(\register_r[23][20] ), .S0(n2556), .S1(n2539), .Y(n2273) );
  MXI4X1 U1477 ( .A(\register_r[20][16] ), .B(\register_r[21][16] ), .C(
        \register_r[22][16] ), .D(\register_r[23][16] ), .S0(n2554), .S1(n2538), .Y(n2241) );
  MXI4X1 U1478 ( .A(\register_r[20][12] ), .B(\register_r[21][12] ), .C(
        \register_r[22][12] ), .D(\register_r[23][12] ), .S0(n2567), .S1(n2546), .Y(n2209) );
  MXI4X1 U1479 ( .A(\register_r[4][12] ), .B(\register_r[5][12] ), .C(
        \register_r[6][12] ), .D(\register_r[7][12] ), .S0(n2565), .S1(n2544), 
        .Y(n2213) );
  MXI4X1 U1480 ( .A(\register_r[20][8] ), .B(\register_r[21][8] ), .C(
        \register_r[22][8] ), .D(\register_r[23][8] ), .S0(n2565), .S1(n2544), 
        .Y(n2177) );
  MXI4X1 U1481 ( .A(\register_r[4][8] ), .B(\register_r[5][8] ), .C(
        \register_r[6][8] ), .D(\register_r[7][8] ), .S0(n2565), .S1(n2544), 
        .Y(n2181) );
  MXI4X1 U1482 ( .A(\register_r[20][4] ), .B(\register_r[21][4] ), .C(
        \register_r[22][4] ), .D(\register_r[23][4] ), .S0(n2563), .S1(n2551), 
        .Y(n2145) );
  MXI4X1 U1483 ( .A(\register_r[4][4] ), .B(\register_r[5][4] ), .C(
        \register_r[6][4] ), .D(\register_r[7][4] ), .S0(n2563), .S1(n2538), 
        .Y(n2149) );
  MXI4X1 U1484 ( .A(\register_r[16][19] ), .B(\register_r[17][19] ), .C(
        \register_r[18][19] ), .D(\register_r[19][19] ), .S0(n3084), .S1(n3066), .Y(n2793) );
  MXI4X1 U1485 ( .A(\register_r[16][18] ), .B(\register_r[17][18] ), .C(
        \register_r[18][18] ), .D(\register_r[19][18] ), .S0(n3084), .S1(n3065), .Y(n2785) );
  MXI4X1 U1486 ( .A(\register_r[16][17] ), .B(\register_r[17][17] ), .C(
        \register_r[18][17] ), .D(\register_r[19][17] ), .S0(n3083), .S1(n3065), .Y(n2777) );
  MXI4X1 U1487 ( .A(\register_r[16][16] ), .B(\register_r[17][16] ), .C(
        \register_r[18][16] ), .D(\register_r[19][16] ), .S0(n3083), .S1(n3065), .Y(n2769) );
  MXI4X1 U1488 ( .A(\register_r[16][31] ), .B(\register_r[17][31] ), .C(
        \register_r[18][31] ), .D(\register_r[19][31] ), .S0(n3090), .S1(n3068), .Y(n2889) );
  MXI4X1 U1489 ( .A(\register_r[16][30] ), .B(\register_r[17][30] ), .C(
        \register_r[18][30] ), .D(\register_r[19][30] ), .S0(n3089), .S1(n3068), .Y(n2881) );
  MXI4X1 U1490 ( .A(\register_r[16][29] ), .B(\register_r[17][29] ), .C(
        \register_r[18][29] ), .D(\register_r[19][29] ), .S0(n3089), .S1(n3068), .Y(n2873) );
  MXI4X1 U1491 ( .A(\register_r[16][28] ), .B(\register_r[17][28] ), .C(
        \register_r[18][28] ), .D(\register_r[19][28] ), .S0(n2559), .S1(n2542), .Y(n2338) );
  MXI4X1 U1492 ( .A(\register_r[16][28] ), .B(\register_r[17][28] ), .C(
        \register_r[18][28] ), .D(\register_r[19][28] ), .S0(n3088), .S1(n3068), .Y(n2865) );
  MXI4X1 U1493 ( .A(\register_r[16][23] ), .B(\register_r[17][23] ), .C(
        \register_r[18][23] ), .D(\register_r[19][23] ), .S0(n3086), .S1(n3072), .Y(n2825) );
  MXI4X1 U1494 ( .A(\register_r[16][22] ), .B(\register_r[17][22] ), .C(
        \register_r[18][22] ), .D(\register_r[19][22] ), .S0(n3086), .S1(n3077), .Y(n2817) );
  MXI4X1 U1495 ( .A(\register_r[16][21] ), .B(\register_r[17][21] ), .C(
        \register_r[18][21] ), .D(\register_r[19][21] ), .S0(n3085), .S1(n3066), .Y(n2809) );
  MXI4X1 U1496 ( .A(\register_r[16][20] ), .B(\register_r[17][20] ), .C(
        \register_r[18][20] ), .D(\register_r[19][20] ), .S0(n3085), .S1(n3066), .Y(n2801) );
  MXI4X1 U1497 ( .A(\register_r[16][26] ), .B(\register_r[17][26] ), .C(
        \register_r[18][26] ), .D(\register_r[19][26] ), .S0(n3087), .S1(n3067), .Y(n2849) );
  MXI4X1 U1498 ( .A(\register_r[16][27] ), .B(\register_r[17][27] ), .C(
        \register_r[18][27] ), .D(\register_r[19][27] ), .S0(n3088), .S1(n3067), .Y(n2857) );
  MXI4X1 U1499 ( .A(\register_r[16][25] ), .B(\register_r[17][25] ), .C(
        \register_r[18][25] ), .D(\register_r[19][25] ), .S0(n3087), .S1(n3067), .Y(n2841) );
  MXI4X1 U1500 ( .A(\register_r[16][24] ), .B(\register_r[17][24] ), .C(
        \register_r[18][24] ), .D(\register_r[19][24] ), .S0(n3087), .S1(n3077), .Y(n2833) );
  MXI4X1 U1501 ( .A(\register_r[16][0] ), .B(\register_r[17][0] ), .C(
        \register_r[18][0] ), .D(\register_r[19][0] ), .S0(n3090), .S1(n3069), 
        .Y(n2641) );
  MXI4X1 U1502 ( .A(\register_r[16][24] ), .B(\register_r[17][24] ), .C(
        \register_r[18][24] ), .D(\register_r[19][24] ), .S0(n2558), .S1(n2540), .Y(n2306) );
  MXI4X1 U1503 ( .A(\register_r[16][20] ), .B(\register_r[17][20] ), .C(
        \register_r[18][20] ), .D(\register_r[19][20] ), .S0(n2556), .S1(n2539), .Y(n2274) );
  MXI4X1 U1504 ( .A(\register_r[16][16] ), .B(\register_r[17][16] ), .C(
        \register_r[18][16] ), .D(\register_r[19][16] ), .S0(n2554), .S1(n2538), .Y(n2242) );
  MXI4X1 U1505 ( .A(\register_r[28][19] ), .B(\register_r[29][19] ), .C(
        \register_r[30][19] ), .D(\register_r[31][19] ), .S0(n3084), .S1(n3065), .Y(n2790) );
  MXI4X1 U1506 ( .A(\register_r[28][18] ), .B(\register_r[29][18] ), .C(
        \register_r[30][18] ), .D(\register_r[31][18] ), .S0(n3083), .S1(n3065), .Y(n2782) );
  MXI4X1 U1507 ( .A(\register_r[28][17] ), .B(\register_r[29][17] ), .C(
        \register_r[30][17] ), .D(\register_r[31][17] ), .S0(n3083), .S1(n3065), .Y(n2774) );
  MXI4X1 U1508 ( .A(\register_r[28][16] ), .B(\register_r[29][16] ), .C(
        \register_r[30][16] ), .D(\register_r[31][16] ), .S0(n3083), .S1(n3065), .Y(n2766) );
  MXI4X1 U1509 ( .A(\register_r[28][31] ), .B(\register_r[29][31] ), .C(
        \register_r[30][31] ), .D(\register_r[31][31] ), .S0(n3090), .S1(n3068), .Y(n2886) );
  MXI4X1 U1510 ( .A(\register_r[28][30] ), .B(\register_r[29][30] ), .C(
        \register_r[30][30] ), .D(\register_r[31][30] ), .S0(n3089), .S1(n3068), .Y(n2878) );
  MXI4X1 U1511 ( .A(\register_r[28][29] ), .B(\register_r[29][29] ), .C(
        \register_r[30][29] ), .D(\register_r[31][29] ), .S0(n3089), .S1(n3068), .Y(n2870) );
  MXI4X1 U1512 ( .A(\register_r[28][28] ), .B(\register_r[29][28] ), .C(
        \register_r[30][28] ), .D(\register_r[31][28] ), .S0(n2559), .S1(n2541), .Y(n2335) );
  MXI4X1 U1513 ( .A(\register_r[28][28] ), .B(\register_r[29][28] ), .C(
        \register_r[30][28] ), .D(\register_r[31][28] ), .S0(n3088), .S1(n3067), .Y(n2862) );
  MXI4X1 U1514 ( .A(\register_r[28][23] ), .B(\register_r[29][23] ), .C(
        \register_r[30][23] ), .D(\register_r[31][23] ), .S0(n3086), .S1(n3069), .Y(n2822) );
  MXI4X1 U1515 ( .A(\register_r[28][22] ), .B(\register_r[29][22] ), .C(
        \register_r[30][22] ), .D(\register_r[31][22] ), .S0(n3085), .S1(n3066), .Y(n2814) );
  MXI4X1 U1516 ( .A(\register_r[28][21] ), .B(\register_r[29][21] ), .C(
        \register_r[30][21] ), .D(\register_r[31][21] ), .S0(n3085), .S1(n3066), .Y(n2806) );
  MXI4X1 U1517 ( .A(\register_r[28][20] ), .B(\register_r[29][20] ), .C(
        \register_r[30][20] ), .D(\register_r[31][20] ), .S0(n3084), .S1(n3066), .Y(n2798) );
  MXI4X1 U1518 ( .A(\register_r[28][26] ), .B(\register_r[29][26] ), .C(
        \register_r[30][26] ), .D(\register_r[31][26] ), .S0(n3087), .S1(n3067), .Y(n2846) );
  MXI4X1 U1519 ( .A(\register_r[28][27] ), .B(\register_r[29][27] ), .C(
        \register_r[30][27] ), .D(\register_r[31][27] ), .S0(n3088), .S1(n3067), .Y(n2854) );
  MXI4X1 U1520 ( .A(\register_r[28][25] ), .B(\register_r[29][25] ), .C(
        \register_r[30][25] ), .D(\register_r[31][25] ), .S0(n3087), .S1(n3078), .Y(n2838) );
  MXI4X1 U1521 ( .A(\register_r[28][24] ), .B(\register_r[29][24] ), .C(
        \register_r[30][24] ), .D(\register_r[31][24] ), .S0(n3086), .S1(n3078), .Y(n2830) );
  MXI4X1 U1522 ( .A(r_12[3]), .B(r_13[3]), .C(\register_r[14][3] ), .D(
        \register_r[15][3] ), .S0(n3081), .S1(n3070), .Y(n2666) );
  MXI4X1 U1523 ( .A(r_12[2]), .B(r_13[2]), .C(\register_r[14][2] ), .D(
        \register_r[15][2] ), .S0(n3091), .S1(n3069), .Y(n2658) );
  MXI4X1 U1524 ( .A(r_12[1]), .B(r_13[1]), .C(\register_r[14][1] ), .D(
        \register_r[15][1] ), .S0(n3091), .S1(n3069), .Y(n2650) );
  MXI4X1 U1525 ( .A(\register_r[28][0] ), .B(\register_r[29][0] ), .C(
        \register_r[30][0] ), .D(\register_r[31][0] ), .S0(n3090), .S1(n3069), 
        .Y(n2638) );
  MXI4X1 U1526 ( .A(r_12[7]), .B(r_13[7]), .C(\register_r[14][7] ), .D(
        \register_r[15][7] ), .S0(n3092), .S1(n3071), .Y(n2698) );
  MXI4X1 U1527 ( .A(r_12[6]), .B(r_13[6]), .C(\register_r[14][6] ), .D(
        \register_r[15][6] ), .S0(n3092), .S1(n3071), .Y(n2690) );
  MXI4X1 U1528 ( .A(r_12[5]), .B(r_13[5]), .C(\register_r[14][5] ), .D(
        \register_r[15][5] ), .S0(n3092), .S1(n3070), .Y(n2682) );
  MXI4X1 U1529 ( .A(r_12[4]), .B(r_13[4]), .C(\register_r[14][4] ), .D(
        \register_r[15][4] ), .S0(n3093), .S1(n3070), .Y(n2674) );
  MXI4X1 U1530 ( .A(r_12[11]), .B(r_13[11]), .C(\register_r[14][11] ), .D(
        \register_r[15][11] ), .S0(n3094), .S1(n3072), .Y(n2730) );
  MXI4X1 U1531 ( .A(r_12[10]), .B(r_13[10]), .C(\register_r[14][10] ), .D(
        \register_r[15][10] ), .S0(n3094), .S1(n3072), .Y(n2722) );
  MXI4X1 U1532 ( .A(r_12[9]), .B(r_13[9]), .C(\register_r[14][9] ), .D(
        \register_r[15][9] ), .S0(n3093), .S1(n3072), .Y(n2714) );
  MXI4X1 U1533 ( .A(r_12[8]), .B(r_13[8]), .C(\register_r[14][8] ), .D(
        \register_r[15][8] ), .S0(n3093), .S1(n3071), .Y(n2706) );
  MXI4X1 U1534 ( .A(r_12[15]), .B(r_13[15]), .C(\register_r[14][15] ), .D(
        \register_r[15][15] ), .S0(n3096), .S1(n3074), .Y(n2762) );
  MXI4X1 U1535 ( .A(r_12[14]), .B(r_13[14]), .C(\register_r[14][14] ), .D(
        \register_r[15][14] ), .S0(n3096), .S1(n3073), .Y(n2754) );
  MXI4X1 U1536 ( .A(r_12[13]), .B(r_13[13]), .C(\register_r[14][13] ), .D(
        \register_r[15][13] ), .S0(n3095), .S1(n3073), .Y(n2746) );
  MXI4X1 U1537 ( .A(r_12[12]), .B(r_13[12]), .C(\register_r[14][12] ), .D(
        \register_r[15][12] ), .S0(n3095), .S1(n3073), .Y(n2738) );
  MXI4X1 U1538 ( .A(\register_r[28][24] ), .B(\register_r[29][24] ), .C(
        \register_r[30][24] ), .D(\register_r[31][24] ), .S0(n2557), .S1(n2540), .Y(n2303) );
  MXI4X1 U1539 ( .A(\register_r[28][20] ), .B(\register_r[29][20] ), .C(
        \register_r[30][20] ), .D(\register_r[31][20] ), .S0(n2555), .S1(n2539), .Y(n2271) );
  MXI4X1 U1540 ( .A(\register_r[28][16] ), .B(\register_r[29][16] ), .C(
        \register_r[30][16] ), .D(\register_r[31][16] ), .S0(n2554), .S1(n2538), .Y(n2239) );
  MXI4X1 U1541 ( .A(r_12[12]), .B(r_13[12]), .C(\register_r[14][12] ), .D(
        \register_r[15][12] ), .S0(n2567), .S1(n2546), .Y(n2211) );
  MXI4X1 U1542 ( .A(r_12[8]), .B(r_13[8]), .C(\register_r[14][8] ), .D(
        \register_r[15][8] ), .S0(n2565), .S1(n2544), .Y(n2179) );
  MXI4X1 U1543 ( .A(r_12[4]), .B(r_13[4]), .C(\register_r[14][4] ), .D(
        \register_r[15][4] ), .S0(n2563), .S1(n2550), .Y(n2147) );
  MXI4X1 U1544 ( .A(\register_r[24][19] ), .B(\register_r[25][19] ), .C(
        \register_r[26][19] ), .D(\register_r[27][19] ), .S0(n3084), .S1(n3066), .Y(n2791) );
  MXI4X1 U1545 ( .A(\register_r[24][18] ), .B(\register_r[25][18] ), .C(
        \register_r[26][18] ), .D(\register_r[27][18] ), .S0(n3084), .S1(n3065), .Y(n2783) );
  MXI4X1 U1546 ( .A(\register_r[24][17] ), .B(\register_r[25][17] ), .C(
        \register_r[26][17] ), .D(\register_r[27][17] ), .S0(n3083), .S1(n3065), .Y(n2775) );
  MXI4X1 U1547 ( .A(\register_r[24][16] ), .B(\register_r[25][16] ), .C(
        \register_r[26][16] ), .D(\register_r[27][16] ), .S0(n3083), .S1(n3065), .Y(n2767) );
  MXI4X1 U1548 ( .A(\register_r[24][31] ), .B(\register_r[25][31] ), .C(
        \register_r[26][31] ), .D(\register_r[27][31] ), .S0(n3090), .S1(n3068), .Y(n2887) );
  MXI4X1 U1549 ( .A(\register_r[24][30] ), .B(\register_r[25][30] ), .C(
        \register_r[26][30] ), .D(\register_r[27][30] ), .S0(n3089), .S1(n3068), .Y(n2879) );
  MXI4X1 U1550 ( .A(\register_r[24][29] ), .B(\register_r[25][29] ), .C(
        \register_r[26][29] ), .D(\register_r[27][29] ), .S0(n3089), .S1(n3068), .Y(n2871) );
  MXI4X1 U1551 ( .A(\register_r[24][28] ), .B(\register_r[25][28] ), .C(
        \register_r[26][28] ), .D(\register_r[27][28] ), .S0(n2559), .S1(n2541), .Y(n2336) );
  MXI4X1 U1552 ( .A(\register_r[24][28] ), .B(\register_r[25][28] ), .C(
        \register_r[26][28] ), .D(\register_r[27][28] ), .S0(n3088), .S1(n3067), .Y(n2863) );
  MXI4X1 U1553 ( .A(\register_r[24][23] ), .B(\register_r[25][23] ), .C(
        \register_r[26][23] ), .D(\register_r[27][23] ), .S0(n3086), .S1(n3069), .Y(n2823) );
  MXI4X1 U1554 ( .A(\register_r[24][22] ), .B(\register_r[25][22] ), .C(
        \register_r[26][22] ), .D(\register_r[27][22] ), .S0(n3085), .S1(n3066), .Y(n2815) );
  MXI4X1 U1555 ( .A(\register_r[24][21] ), .B(\register_r[25][21] ), .C(
        \register_r[26][21] ), .D(\register_r[27][21] ), .S0(n3085), .S1(n3066), .Y(n2807) );
  MXI4X1 U1556 ( .A(\register_r[24][20] ), .B(\register_r[25][20] ), .C(
        \register_r[26][20] ), .D(\register_r[27][20] ), .S0(n3084), .S1(n3066), .Y(n2799) );
  MXI4X1 U1557 ( .A(\register_r[24][26] ), .B(\register_r[25][26] ), .C(
        \register_r[26][26] ), .D(\register_r[27][26] ), .S0(n3087), .S1(n3067), .Y(n2847) );
  MXI4X1 U1558 ( .A(\register_r[24][27] ), .B(\register_r[25][27] ), .C(
        \register_r[26][27] ), .D(\register_r[27][27] ), .S0(n3088), .S1(n3067), .Y(n2855) );
  MXI4X1 U1559 ( .A(\register_r[24][25] ), .B(\register_r[25][25] ), .C(
        \register_r[26][25] ), .D(\register_r[27][25] ), .S0(n3087), .S1(n3077), .Y(n2839) );
  MXI4X1 U1560 ( .A(\register_r[24][24] ), .B(\register_r[25][24] ), .C(
        \register_r[26][24] ), .D(\register_r[27][24] ), .S0(n3086), .S1(n3078), .Y(n2831) );
  MXI4X1 U1561 ( .A(\register_r[8][3] ), .B(\register_r[9][3] ), .C(
        \register_r[10][3] ), .D(\register_r[11][3] ), .S0(n3081), .S1(n3070), 
        .Y(n2667) );
  MXI4X1 U1562 ( .A(\register_r[8][2] ), .B(\register_r[9][2] ), .C(
        \register_r[10][2] ), .D(\register_r[11][2] ), .S0(n3091), .S1(n3069), 
        .Y(n2659) );
  MXI4X1 U1563 ( .A(\register_r[8][1] ), .B(\register_r[9][1] ), .C(
        \register_r[10][1] ), .D(\register_r[11][1] ), .S0(n3091), .S1(n3069), 
        .Y(n2651) );
  MXI4X1 U1564 ( .A(\register_r[24][0] ), .B(\register_r[25][0] ), .C(
        \register_r[26][0] ), .D(\register_r[27][0] ), .S0(n3090), .S1(n3069), 
        .Y(n2639) );
  MXI4X1 U1565 ( .A(\register_r[8][7] ), .B(\register_r[9][7] ), .C(
        \register_r[10][7] ), .D(\register_r[11][7] ), .S0(n3093), .S1(n3071), 
        .Y(n2699) );
  MXI4X1 U1566 ( .A(\register_r[8][6] ), .B(\register_r[9][6] ), .C(
        \register_r[10][6] ), .D(\register_r[11][6] ), .S0(n3092), .S1(n3071), 
        .Y(n2691) );
  MXI4X1 U1567 ( .A(\register_r[8][5] ), .B(\register_r[9][5] ), .C(
        \register_r[10][5] ), .D(\register_r[11][5] ), .S0(n3092), .S1(n3070), 
        .Y(n2683) );
  MXI4X1 U1568 ( .A(\register_r[8][4] ), .B(\register_r[9][4] ), .C(
        \register_r[10][4] ), .D(\register_r[11][4] ), .S0(n3081), .S1(n3070), 
        .Y(n2675) );
  MXI4X1 U1569 ( .A(\register_r[8][11] ), .B(\register_r[9][11] ), .C(
        \register_r[10][11] ), .D(\register_r[11][11] ), .S0(n3094), .S1(n3072), .Y(n2731) );
  MXI4X1 U1570 ( .A(\register_r[8][10] ), .B(\register_r[9][10] ), .C(
        \register_r[10][10] ), .D(\register_r[11][10] ), .S0(n3094), .S1(n3072), .Y(n2723) );
  MXI4X1 U1571 ( .A(\register_r[8][9] ), .B(\register_r[9][9] ), .C(
        \register_r[10][9] ), .D(\register_r[11][9] ), .S0(n3094), .S1(n3072), 
        .Y(n2715) );
  MXI4X1 U1572 ( .A(\register_r[8][8] ), .B(\register_r[9][8] ), .C(
        \register_r[10][8] ), .D(\register_r[11][8] ), .S0(n3093), .S1(n3071), 
        .Y(n2707) );
  MXI4X1 U1573 ( .A(\register_r[8][15] ), .B(\register_r[9][15] ), .C(
        \register_r[10][15] ), .D(\register_r[11][15] ), .S0(n3096), .S1(n3074), .Y(n2763) );
  MXI4X1 U1574 ( .A(\register_r[8][14] ), .B(\register_r[9][14] ), .C(
        \register_r[10][14] ), .D(\register_r[11][14] ), .S0(n3096), .S1(n3073), .Y(n2755) );
  MXI4X1 U1575 ( .A(\register_r[8][13] ), .B(\register_r[9][13] ), .C(
        \register_r[10][13] ), .D(\register_r[11][13] ), .S0(n3095), .S1(n3073), .Y(n2747) );
  MXI4X1 U1576 ( .A(\register_r[8][12] ), .B(\register_r[9][12] ), .C(
        \register_r[10][12] ), .D(\register_r[11][12] ), .S0(n3095), .S1(n3073), .Y(n2739) );
  MXI4X1 U1577 ( .A(\register_r[24][24] ), .B(\register_r[25][24] ), .C(
        \register_r[26][24] ), .D(\register_r[27][24] ), .S0(n2557), .S1(n2540), .Y(n2304) );
  MXI4X1 U1578 ( .A(\register_r[24][20] ), .B(\register_r[25][20] ), .C(
        \register_r[26][20] ), .D(\register_r[27][20] ), .S0(n2555), .S1(n2539), .Y(n2272) );
  MXI4X1 U1579 ( .A(\register_r[24][16] ), .B(\register_r[25][16] ), .C(
        \register_r[26][16] ), .D(\register_r[27][16] ), .S0(n2554), .S1(n2538), .Y(n2240) );
  MXI4X1 U1580 ( .A(\register_r[8][12] ), .B(\register_r[9][12] ), .C(
        \register_r[10][12] ), .D(\register_r[11][12] ), .S0(n2567), .S1(n2546), .Y(n2212) );
  MXI4X1 U1581 ( .A(\register_r[8][8] ), .B(\register_r[9][8] ), .C(
        \register_r[10][8] ), .D(\register_r[11][8] ), .S0(n2565), .S1(n2544), 
        .Y(n2180) );
  MXI4X1 U1582 ( .A(\register_r[8][4] ), .B(\register_r[9][4] ), .C(
        \register_r[10][4] ), .D(\register_r[11][4] ), .S0(n2563), .S1(n2538), 
        .Y(n2148) );
  NOR2X2 U1583 ( .A(WriteReg[1]), .B(WriteReg[2]), .Y(n43) );
  NOR2BX1 U1584 ( .AN(n59), .B(WriteReg[0]), .Y(n48) );
  CLKINVX1 U1585 ( .A(WriteReg[0]), .Y(n3441) );
  NOR3X1 U1586 ( .A(WriteReg[3]), .B(WriteReg[4]), .C(n3440), .Y(n59) );
  NOR3X1 U1587 ( .A(n3440), .B(WriteReg[4]), .C(n3442), .Y(n80) );
  CLKINVX1 U1588 ( .A(WriteReg[1]), .Y(n3444) );
  OAI22XL U1589 ( .A0(n3165), .A1(n3291), .B0(n3289), .B1(n1098), .Y(n1163) );
  OAI22XL U1590 ( .A0(n3163), .A1(n3291), .B0(n3289), .B1(n1097), .Y(n1164) );
  OAI22XL U1591 ( .A0(n3161), .A1(n3291), .B0(n3289), .B1(n1096), .Y(n1165) );
  OAI22XL U1592 ( .A0(n3159), .A1(n3291), .B0(n3289), .B1(n1095), .Y(n1166) );
  OAI22XL U1593 ( .A0(n3157), .A1(n3288), .B0(n3289), .B1(n1094), .Y(n1167) );
  OAI22XL U1594 ( .A0(n3155), .A1(n3288), .B0(n3289), .B1(n1093), .Y(n1168) );
  OAI22XL U1595 ( .A0(n3153), .A1(n3288), .B0(n3289), .B1(n1092), .Y(n1169) );
  OAI22XL U1596 ( .A0(n3151), .A1(n3288), .B0(n3289), .B1(n1091), .Y(n1170) );
  OAI22XL U1597 ( .A0(n3149), .A1(n3288), .B0(n3289), .B1(n1090), .Y(n1171) );
  OAI22XL U1598 ( .A0(n3147), .A1(n3288), .B0(n3289), .B1(n1089), .Y(n1172) );
  OAI22XL U1599 ( .A0(n3145), .A1(n3291), .B0(n3289), .B1(n1088), .Y(n1173) );
  OAI22XL U1600 ( .A0(n3143), .A1(n3291), .B0(n3289), .B1(n1087), .Y(n1174) );
  OAI22XL U1601 ( .A0(n3141), .A1(n45), .B0(n3290), .B1(n1086), .Y(n1175) );
  OAI22XL U1602 ( .A0(n3139), .A1(n3288), .B0(n3290), .B1(n1085), .Y(n1176) );
  OAI22XL U1603 ( .A0(n3137), .A1(n3288), .B0(n3290), .B1(n1084), .Y(n1177) );
  OAI22XL U1604 ( .A0(n3135), .A1(n3288), .B0(n3290), .B1(n1083), .Y(n1178) );
  OAI22XL U1605 ( .A0(n3133), .A1(n3288), .B0(n3289), .B1(n1082), .Y(n1179) );
  OAI22XL U1606 ( .A0(n3131), .A1(n3288), .B0(n3290), .B1(n1081), .Y(n1180) );
  OAI22XL U1607 ( .A0(n3129), .A1(n45), .B0(n3289), .B1(n1080), .Y(n1181) );
  OAI22XL U1608 ( .A0(n3127), .A1(n45), .B0(n3290), .B1(n1079), .Y(n1182) );
  OAI22XL U1609 ( .A0(n3125), .A1(n3291), .B0(n3289), .B1(n1078), .Y(n1183) );
  OAI22XL U1610 ( .A0(n3123), .A1(n3288), .B0(n3290), .B1(n1077), .Y(n1184) );
  OAI22XL U1611 ( .A0(n3121), .A1(n3291), .B0(n3289), .B1(n1076), .Y(n1185) );
  OAI22XL U1612 ( .A0(n3119), .A1(n3288), .B0(n3290), .B1(n1075), .Y(n1186) );
  OAI22XL U1613 ( .A0(n3117), .A1(n45), .B0(n3290), .B1(n1074), .Y(n1187) );
  OAI22XL U1614 ( .A0(n3115), .A1(n3291), .B0(n3290), .B1(n1073), .Y(n1188) );
  OAI22XL U1615 ( .A0(n3113), .A1(n3288), .B0(n3290), .B1(n1072), .Y(n1189) );
  OAI22XL U1616 ( .A0(n3111), .A1(n3288), .B0(n3290), .B1(n1071), .Y(n1190) );
  OAI22XL U1617 ( .A0(n3109), .A1(n3288), .B0(n3290), .B1(n1070), .Y(n1191) );
  OAI22XL U1618 ( .A0(n3107), .A1(n3288), .B0(n3290), .B1(n1069), .Y(n1192) );
  OAI22XL U1619 ( .A0(n3105), .A1(n3288), .B0(n3290), .B1(n1068), .Y(n1193) );
  OAI22XL U1620 ( .A0(n3103), .A1(n3291), .B0(n3290), .B1(n1067), .Y(n1194) );
  OAI22XL U1621 ( .A0(n3165), .A1(n3287), .B0(n3285), .B1(n1066), .Y(n1195) );
  OAI22XL U1622 ( .A0(n3163), .A1(n3287), .B0(n3285), .B1(n1065), .Y(n1196) );
  OAI22XL U1623 ( .A0(n3161), .A1(n3287), .B0(n3285), .B1(n1064), .Y(n1197) );
  OAI22XL U1624 ( .A0(n3159), .A1(n3287), .B0(n3285), .B1(n1063), .Y(n1198) );
  OAI22XL U1625 ( .A0(n3157), .A1(n3284), .B0(n3285), .B1(n1062), .Y(n1199) );
  OAI22XL U1626 ( .A0(n3155), .A1(n3284), .B0(n3285), .B1(n1061), .Y(n1200) );
  OAI22XL U1627 ( .A0(n3153), .A1(n3284), .B0(n3285), .B1(n1060), .Y(n1201) );
  OAI22XL U1628 ( .A0(n3151), .A1(n49), .B0(n3285), .B1(n1059), .Y(n1202) );
  OAI22XL U1629 ( .A0(n3149), .A1(n3287), .B0(n3285), .B1(n1058), .Y(n1203) );
  OAI22XL U1630 ( .A0(n3147), .A1(n3287), .B0(n3285), .B1(n1057), .Y(n1204) );
  OAI22XL U1631 ( .A0(n3145), .A1(n3287), .B0(n3285), .B1(n1056), .Y(n1205) );
  OAI22XL U1632 ( .A0(n3143), .A1(n3287), .B0(n3285), .B1(n1055), .Y(n1206) );
  OAI22XL U1633 ( .A0(n3141), .A1(n3284), .B0(n3286), .B1(n1054), .Y(n1207) );
  OAI22XL U1634 ( .A0(n3139), .A1(n3284), .B0(n3286), .B1(n1053), .Y(n1208) );
  OAI22XL U1635 ( .A0(n3137), .A1(n3284), .B0(n3286), .B1(n1052), .Y(n1209) );
  OAI22XL U1636 ( .A0(n3135), .A1(n3284), .B0(n3286), .B1(n1051), .Y(n1210) );
  OAI22XL U1637 ( .A0(n3133), .A1(n49), .B0(n3285), .B1(n1050), .Y(n1211) );
  OAI22XL U1638 ( .A0(n3131), .A1(n49), .B0(n3286), .B1(n1049), .Y(n1212) );
  OAI22XL U1639 ( .A0(n3129), .A1(n49), .B0(n3285), .B1(n1048), .Y(n1213) );
  OAI22XL U1640 ( .A0(n3127), .A1(n3284), .B0(n3286), .B1(n1047), .Y(n1214) );
  OAI22XL U1641 ( .A0(n3125), .A1(n3287), .B0(n3285), .B1(n1046), .Y(n1215) );
  OAI22XL U1642 ( .A0(n3123), .A1(n3284), .B0(n3286), .B1(n1045), .Y(n1216) );
  OAI22XL U1643 ( .A0(n3121), .A1(n3284), .B0(n3285), .B1(n1044), .Y(n1217) );
  OAI22XL U1644 ( .A0(n3119), .A1(n3284), .B0(n3286), .B1(n1043), .Y(n1218) );
  OAI22XL U1645 ( .A0(n3165), .A1(n3283), .B0(n3281), .B1(n1034), .Y(n1227) );
  OAI22XL U1646 ( .A0(n3163), .A1(n3283), .B0(n3281), .B1(n1033), .Y(n1228) );
  OAI22XL U1647 ( .A0(n3161), .A1(n3283), .B0(n3281), .B1(n1032), .Y(n1229) );
  OAI22XL U1648 ( .A0(n3159), .A1(n3283), .B0(n3281), .B1(n1031), .Y(n1230) );
  OAI22XL U1649 ( .A0(n3157), .A1(n3283), .B0(n3281), .B1(n1030), .Y(n1231) );
  OAI22XL U1650 ( .A0(n3155), .A1(n3283), .B0(n3281), .B1(n1029), .Y(n1232) );
  OAI22XL U1651 ( .A0(n3153), .A1(n3283), .B0(n3281), .B1(n1028), .Y(n1233) );
  OAI22XL U1652 ( .A0(n3151), .A1(n3283), .B0(n3281), .B1(n1027), .Y(n1234) );
  OAI22XL U1653 ( .A0(n3149), .A1(n3283), .B0(n3281), .B1(n1026), .Y(n1235) );
  OAI22XL U1654 ( .A0(n3147), .A1(n3283), .B0(n3281), .B1(n1025), .Y(n1236) );
  OAI22XL U1655 ( .A0(n3145), .A1(n3283), .B0(n3281), .B1(n1024), .Y(n1237) );
  OAI22XL U1656 ( .A0(n3143), .A1(n3283), .B0(n3281), .B1(n1023), .Y(n1238) );
  OAI22XL U1657 ( .A0(n3141), .A1(n3280), .B0(n3282), .B1(n1022), .Y(n1239) );
  OAI22XL U1658 ( .A0(n3139), .A1(n3280), .B0(n3282), .B1(n1021), .Y(n1240) );
  OAI22XL U1659 ( .A0(n3137), .A1(n3280), .B0(n3282), .B1(n1020), .Y(n1241) );
  OAI22XL U1660 ( .A0(n3135), .A1(n3280), .B0(n3282), .B1(n1019), .Y(n1242) );
  OAI22XL U1661 ( .A0(n3133), .A1(n3280), .B0(n3282), .B1(n1018), .Y(n1243) );
  OAI22XL U1662 ( .A0(n3131), .A1(n3283), .B0(n3282), .B1(n1017), .Y(n1244) );
  OAI22XL U1663 ( .A0(n3129), .A1(n3283), .B0(n3282), .B1(n1016), .Y(n1245) );
  OAI22XL U1664 ( .A0(n3127), .A1(n3280), .B0(n3282), .B1(n1015), .Y(n1246) );
  OAI22XL U1665 ( .A0(n3125), .A1(n3280), .B0(n3282), .B1(n1014), .Y(n1247) );
  OAI22XL U1666 ( .A0(n3123), .A1(n3283), .B0(n3282), .B1(n1013), .Y(n1248) );
  OAI22XL U1667 ( .A0(n3121), .A1(n3280), .B0(n3282), .B1(n1012), .Y(n1249) );
  OAI22XL U1668 ( .A0(n3119), .A1(n3283), .B0(n3282), .B1(n1011), .Y(n1250) );
  OAI22XL U1669 ( .A0(n3165), .A1(n3279), .B0(n3277), .B1(n1002), .Y(n1259) );
  OAI22XL U1670 ( .A0(n3163), .A1(n3279), .B0(n3277), .B1(n1001), .Y(n1260) );
  OAI22XL U1671 ( .A0(n3161), .A1(n3279), .B0(n3277), .B1(n1000), .Y(n1261) );
  OAI22XL U1672 ( .A0(n3159), .A1(n3279), .B0(n3277), .B1(n999), .Y(n1262) );
  OAI22XL U1673 ( .A0(n3157), .A1(n3276), .B0(n3277), .B1(n998), .Y(n1263) );
  OAI22XL U1674 ( .A0(n3155), .A1(n3276), .B0(n3277), .B1(n997), .Y(n1264) );
  OAI22XL U1675 ( .A0(n3153), .A1(n3276), .B0(n3277), .B1(n996), .Y(n1265) );
  OAI22XL U1676 ( .A0(n3151), .A1(n54), .B0(n3277), .B1(n995), .Y(n1266) );
  OAI22XL U1677 ( .A0(n3149), .A1(n3279), .B0(n3277), .B1(n994), .Y(n1267) );
  OAI22XL U1678 ( .A0(n3147), .A1(n3279), .B0(n3277), .B1(n993), .Y(n1268) );
  OAI22XL U1679 ( .A0(n3145), .A1(n3279), .B0(n3277), .B1(n992), .Y(n1269) );
  OAI22XL U1680 ( .A0(n3143), .A1(n3279), .B0(n3277), .B1(n991), .Y(n1270) );
  OAI22XL U1681 ( .A0(n3141), .A1(n3276), .B0(n3278), .B1(n990), .Y(n1271) );
  OAI22XL U1682 ( .A0(n3139), .A1(n3276), .B0(n3278), .B1(n989), .Y(n1272) );
  OAI22XL U1683 ( .A0(n3137), .A1(n3276), .B0(n3278), .B1(n988), .Y(n1273) );
  OAI22XL U1684 ( .A0(n3135), .A1(n3276), .B0(n3278), .B1(n987), .Y(n1274) );
  OAI22XL U1685 ( .A0(n3133), .A1(n54), .B0(n3278), .B1(n986), .Y(n1275) );
  OAI22XL U1686 ( .A0(n3131), .A1(n54), .B0(n3278), .B1(n985), .Y(n1276) );
  OAI22XL U1687 ( .A0(n3129), .A1(n54), .B0(n3278), .B1(n984), .Y(n1277) );
  OAI22XL U1688 ( .A0(n3127), .A1(n3276), .B0(n3278), .B1(n983), .Y(n1278) );
  OAI22XL U1689 ( .A0(n3125), .A1(n3279), .B0(n3278), .B1(n982), .Y(n1279) );
  OAI22XL U1690 ( .A0(n3123), .A1(n3276), .B0(n3278), .B1(n981), .Y(n1280) );
  OAI22XL U1691 ( .A0(n3121), .A1(n3276), .B0(n3278), .B1(n980), .Y(n1281) );
  OAI22XL U1692 ( .A0(n3119), .A1(n3276), .B0(n3278), .B1(n979), .Y(n1282) );
  OAI22XL U1693 ( .A0(n3165), .A1(n3275), .B0(n3273), .B1(n970), .Y(n1291) );
  OAI22XL U1694 ( .A0(n3163), .A1(n3275), .B0(n3273), .B1(n969), .Y(n1292) );
  OAI22XL U1695 ( .A0(n3161), .A1(n3275), .B0(n3273), .B1(n968), .Y(n1293) );
  OAI22XL U1696 ( .A0(n3159), .A1(n3275), .B0(n3273), .B1(n967), .Y(n1294) );
  OAI22XL U1697 ( .A0(n3157), .A1(n3275), .B0(n3273), .B1(n966), .Y(n1295) );
  OAI22XL U1698 ( .A0(n3155), .A1(n3275), .B0(n3273), .B1(n965), .Y(n1296) );
  OAI22XL U1699 ( .A0(n3153), .A1(n3275), .B0(n3273), .B1(n964), .Y(n1297) );
  OAI22XL U1700 ( .A0(n3151), .A1(n3275), .B0(n3273), .B1(n963), .Y(n1298) );
  OAI22XL U1701 ( .A0(n3149), .A1(n3275), .B0(n3273), .B1(n962), .Y(n1299) );
  OAI22XL U1702 ( .A0(n3147), .A1(n3275), .B0(n3273), .B1(n961), .Y(n1300) );
  OAI22XL U1703 ( .A0(n3145), .A1(n3275), .B0(n3273), .B1(n960), .Y(n1301) );
  OAI22XL U1704 ( .A0(n3143), .A1(n3275), .B0(n3273), .B1(n959), .Y(n1302) );
  OAI22XL U1705 ( .A0(n3141), .A1(n3272), .B0(n3274), .B1(n958), .Y(n1303) );
  OAI22XL U1706 ( .A0(n3139), .A1(n3272), .B0(n3274), .B1(n957), .Y(n1304) );
  OAI22XL U1707 ( .A0(n3137), .A1(n3272), .B0(n3274), .B1(n956), .Y(n1305) );
  OAI22XL U1708 ( .A0(n3135), .A1(n3272), .B0(n3274), .B1(n955), .Y(n1306) );
  OAI22XL U1709 ( .A0(n3133), .A1(n3272), .B0(n3274), .B1(n954), .Y(n1307) );
  OAI22XL U1710 ( .A0(n3131), .A1(n3275), .B0(n3274), .B1(n953), .Y(n1308) );
  OAI22XL U1711 ( .A0(n3129), .A1(n3275), .B0(n3274), .B1(n952), .Y(n1309) );
  OAI22XL U1712 ( .A0(n3127), .A1(n3272), .B0(n3274), .B1(n951), .Y(n1310) );
  OAI22XL U1713 ( .A0(n3125), .A1(n3272), .B0(n3274), .B1(n950), .Y(n1311) );
  OAI22XL U1714 ( .A0(n3123), .A1(n3275), .B0(n3274), .B1(n949), .Y(n1312) );
  OAI22XL U1715 ( .A0(n3121), .A1(n3272), .B0(n3274), .B1(n948), .Y(n1313) );
  OAI22XL U1716 ( .A0(n3119), .A1(n3275), .B0(n3274), .B1(n947), .Y(n1314) );
  OAI22XL U1717 ( .A0(n3165), .A1(n3271), .B0(n3269), .B1(n938), .Y(n1323) );
  OAI22XL U1718 ( .A0(n3163), .A1(n3271), .B0(n3269), .B1(n937), .Y(n1324) );
  OAI22XL U1719 ( .A0(n3161), .A1(n3271), .B0(n3269), .B1(n936), .Y(n1325) );
  OAI22XL U1720 ( .A0(n3159), .A1(n3271), .B0(n3269), .B1(n935), .Y(n1326) );
  OAI22XL U1721 ( .A0(n3157), .A1(n3268), .B0(n3269), .B1(n934), .Y(n1327) );
  OAI22XL U1722 ( .A0(n3155), .A1(n3268), .B0(n3269), .B1(n933), .Y(n1328) );
  OAI22XL U1723 ( .A0(n3153), .A1(n3268), .B0(n3269), .B1(n932), .Y(n1329) );
  OAI22XL U1724 ( .A0(n3151), .A1(n60), .B0(n3269), .B1(n931), .Y(n1330) );
  OAI22XL U1725 ( .A0(n3149), .A1(n3271), .B0(n3269), .B1(n930), .Y(n1331) );
  OAI22XL U1726 ( .A0(n3147), .A1(n3271), .B0(n3269), .B1(n929), .Y(n1332) );
  OAI22XL U1727 ( .A0(n3145), .A1(n3271), .B0(n3269), .B1(n928), .Y(n1333) );
  OAI22XL U1728 ( .A0(n3143), .A1(n3271), .B0(n3269), .B1(n927), .Y(n1334) );
  OAI22XL U1729 ( .A0(n3141), .A1(n3268), .B0(n3270), .B1(n926), .Y(n1335) );
  OAI22XL U1730 ( .A0(n3139), .A1(n3268), .B0(n3270), .B1(n925), .Y(n1336) );
  OAI22XL U1731 ( .A0(n3137), .A1(n3268), .B0(n3270), .B1(n924), .Y(n1337) );
  OAI22XL U1732 ( .A0(n3135), .A1(n3268), .B0(n3270), .B1(n923), .Y(n1338) );
  OAI22XL U1733 ( .A0(n3133), .A1(n60), .B0(n3270), .B1(n922), .Y(n1339) );
  OAI22XL U1734 ( .A0(n3131), .A1(n60), .B0(n3270), .B1(n921), .Y(n1340) );
  OAI22XL U1735 ( .A0(n3129), .A1(n60), .B0(n3270), .B1(n920), .Y(n1341) );
  OAI22XL U1736 ( .A0(n3127), .A1(n3268), .B0(n3270), .B1(n919), .Y(n1342) );
  OAI22XL U1737 ( .A0(n3125), .A1(n3271), .B0(n3270), .B1(n918), .Y(n1343) );
  OAI22XL U1738 ( .A0(n3123), .A1(n3268), .B0(n3270), .B1(n917), .Y(n1344) );
  OAI22XL U1739 ( .A0(n3121), .A1(n3268), .B0(n3270), .B1(n916), .Y(n1345) );
  OAI22XL U1740 ( .A0(n3119), .A1(n3268), .B0(n3270), .B1(n915), .Y(n1346) );
  OAI22XL U1741 ( .A0(n3165), .A1(n3267), .B0(n3265), .B1(n906), .Y(n1355) );
  OAI22XL U1742 ( .A0(n3163), .A1(n3267), .B0(n3265), .B1(n905), .Y(n1356) );
  OAI22XL U1743 ( .A0(n3161), .A1(n3267), .B0(n3265), .B1(n904), .Y(n1357) );
  OAI22XL U1744 ( .A0(n3159), .A1(n3267), .B0(n3265), .B1(n903), .Y(n1358) );
  OAI22XL U1745 ( .A0(n3157), .A1(n3264), .B0(n3265), .B1(n902), .Y(n1359) );
  OAI22XL U1746 ( .A0(n3155), .A1(n3267), .B0(n3265), .B1(n901), .Y(n1360) );
  OAI22XL U1747 ( .A0(n3153), .A1(n3264), .B0(n3265), .B1(n900), .Y(n1361) );
  OAI22XL U1748 ( .A0(n3151), .A1(n3264), .B0(n3265), .B1(n899), .Y(n1362) );
  OAI22XL U1749 ( .A0(n3149), .A1(n3267), .B0(n3265), .B1(n898), .Y(n1363) );
  OAI22XL U1750 ( .A0(n3147), .A1(n3267), .B0(n3265), .B1(n897), .Y(n1364) );
  OAI22XL U1751 ( .A0(n3145), .A1(n3264), .B0(n3265), .B1(n896), .Y(n1365) );
  OAI22XL U1752 ( .A0(n3143), .A1(n3267), .B0(n3265), .B1(n895), .Y(n1366) );
  OAI22XL U1753 ( .A0(n3141), .A1(n3264), .B0(n3266), .B1(n894), .Y(n1367) );
  OAI22XL U1754 ( .A0(n3139), .A1(n3264), .B0(n3266), .B1(n893), .Y(n1368) );
  OAI22XL U1755 ( .A0(n3137), .A1(n3264), .B0(n3266), .B1(n892), .Y(n1369) );
  OAI22XL U1756 ( .A0(n3135), .A1(n3264), .B0(n3266), .B1(n891), .Y(n1370) );
  OAI22XL U1757 ( .A0(n3133), .A1(n64), .B0(n3266), .B1(n890), .Y(n1371) );
  OAI22XL U1758 ( .A0(n3131), .A1(n64), .B0(n3266), .B1(n889), .Y(n1372) );
  OAI22XL U1759 ( .A0(n3129), .A1(n64), .B0(n3266), .B1(n888), .Y(n1373) );
  OAI22XL U1760 ( .A0(n3127), .A1(n64), .B0(n3266), .B1(n887), .Y(n1374) );
  OAI22XL U1761 ( .A0(n3125), .A1(n64), .B0(n3266), .B1(n886), .Y(n1375) );
  OAI22XL U1762 ( .A0(n3123), .A1(n3264), .B0(n3266), .B1(n885), .Y(n1376) );
  OAI22XL U1763 ( .A0(n3121), .A1(n3264), .B0(n3266), .B1(n884), .Y(n1377) );
  OAI22XL U1764 ( .A0(n3119), .A1(n3264), .B0(n3266), .B1(n883), .Y(n1378) );
  OAI22XL U1765 ( .A0(n3165), .A1(n3263), .B0(n3261), .B1(n874), .Y(n1387) );
  OAI22XL U1766 ( .A0(n3163), .A1(n3263), .B0(n3261), .B1(n873), .Y(n1388) );
  OAI22XL U1767 ( .A0(n3161), .A1(n3263), .B0(n3261), .B1(n872), .Y(n1389) );
  OAI22XL U1768 ( .A0(n3159), .A1(n3263), .B0(n3261), .B1(n871), .Y(n1390) );
  OAI22XL U1769 ( .A0(n3157), .A1(n3260), .B0(n3261), .B1(n870), .Y(n1391) );
  OAI22XL U1770 ( .A0(n3155), .A1(n3263), .B0(n3261), .B1(n869), .Y(n1392) );
  OAI22XL U1771 ( .A0(n3153), .A1(n3260), .B0(n3261), .B1(n868), .Y(n1393) );
  OAI22XL U1772 ( .A0(n3151), .A1(n3260), .B0(n3261), .B1(n867), .Y(n1394) );
  OAI22XL U1773 ( .A0(n3149), .A1(n3263), .B0(n3261), .B1(n866), .Y(n1395) );
  OAI22XL U1774 ( .A0(n3147), .A1(n3263), .B0(n3261), .B1(n865), .Y(n1396) );
  OAI22XL U1775 ( .A0(n3145), .A1(n3260), .B0(n3261), .B1(n864), .Y(n1397) );
  OAI22XL U1776 ( .A0(n3143), .A1(n3263), .B0(n3261), .B1(n863), .Y(n1398) );
  OAI22XL U1777 ( .A0(n3141), .A1(n3260), .B0(n3262), .B1(n862), .Y(n1399) );
  OAI22XL U1778 ( .A0(n3139), .A1(n3260), .B0(n3262), .B1(n861), .Y(n1400) );
  OAI22XL U1779 ( .A0(n3137), .A1(n3260), .B0(n3262), .B1(n860), .Y(n1401) );
  OAI22XL U1780 ( .A0(n3135), .A1(n3260), .B0(n3262), .B1(n859), .Y(n1402) );
  OAI22XL U1781 ( .A0(n3133), .A1(n67), .B0(n3262), .B1(n858), .Y(n1403) );
  OAI22XL U1782 ( .A0(n3131), .A1(n67), .B0(n3262), .B1(n857), .Y(n1404) );
  OAI22XL U1783 ( .A0(n3129), .A1(n67), .B0(n3262), .B1(n856), .Y(n1405) );
  OAI22XL U1784 ( .A0(n3127), .A1(n67), .B0(n3262), .B1(n855), .Y(n1406) );
  OAI22XL U1785 ( .A0(n3125), .A1(n67), .B0(n3262), .B1(n854), .Y(n1407) );
  OAI22XL U1786 ( .A0(n3123), .A1(n3260), .B0(n3262), .B1(n853), .Y(n1408) );
  OAI22XL U1787 ( .A0(n3121), .A1(n3260), .B0(n3262), .B1(n852), .Y(n1409) );
  OAI22XL U1788 ( .A0(n3119), .A1(n3260), .B0(n3262), .B1(n851), .Y(n1410) );
  OAI22XL U1789 ( .A0(n3165), .A1(n3259), .B0(n3257), .B1(n842), .Y(n1419) );
  OAI22XL U1790 ( .A0(n3163), .A1(n3259), .B0(n3257), .B1(n841), .Y(n1420) );
  OAI22XL U1791 ( .A0(n3161), .A1(n3259), .B0(n3257), .B1(n840), .Y(n1421) );
  OAI22XL U1792 ( .A0(n3159), .A1(n3259), .B0(n3257), .B1(n839), .Y(n1422) );
  OAI22XL U1793 ( .A0(n3157), .A1(n3256), .B0(n3257), .B1(n838), .Y(n1423) );
  OAI22XL U1794 ( .A0(n3155), .A1(n3259), .B0(n3257), .B1(n837), .Y(n1424) );
  OAI22XL U1795 ( .A0(n3153), .A1(n3256), .B0(n3257), .B1(n836), .Y(n1425) );
  OAI22XL U1796 ( .A0(n3151), .A1(n3256), .B0(n3257), .B1(n835), .Y(n1426) );
  OAI22XL U1797 ( .A0(n3149), .A1(n3259), .B0(n3257), .B1(n834), .Y(n1427) );
  OAI22XL U1798 ( .A0(n3147), .A1(n3259), .B0(n3257), .B1(n833), .Y(n1428) );
  OAI22XL U1799 ( .A0(n3145), .A1(n3256), .B0(n3257), .B1(n832), .Y(n1429) );
  OAI22XL U1800 ( .A0(n3143), .A1(n3259), .B0(n3257), .B1(n831), .Y(n1430) );
  OAI22XL U1801 ( .A0(n3141), .A1(n3256), .B0(n3258), .B1(n830), .Y(n1431) );
  OAI22XL U1802 ( .A0(n3139), .A1(n3256), .B0(n3258), .B1(n829), .Y(n1432) );
  OAI22XL U1803 ( .A0(n3137), .A1(n3256), .B0(n3258), .B1(n828), .Y(n1433) );
  OAI22XL U1804 ( .A0(n3135), .A1(n3256), .B0(n3258), .B1(n827), .Y(n1434) );
  OAI22XL U1805 ( .A0(n3133), .A1(n70), .B0(n3258), .B1(n826), .Y(n1435) );
  OAI22XL U1806 ( .A0(n3131), .A1(n70), .B0(n3258), .B1(n825), .Y(n1436) );
  OAI22XL U1807 ( .A0(n3129), .A1(n70), .B0(n3258), .B1(n824), .Y(n1437) );
  OAI22XL U1808 ( .A0(n3127), .A1(n70), .B0(n3258), .B1(n823), .Y(n1438) );
  OAI22XL U1809 ( .A0(n3125), .A1(n70), .B0(n3258), .B1(n822), .Y(n1439) );
  OAI22XL U1810 ( .A0(n3123), .A1(n3256), .B0(n3258), .B1(n821), .Y(n1440) );
  OAI22XL U1811 ( .A0(n3121), .A1(n3256), .B0(n3258), .B1(n820), .Y(n1441) );
  OAI22XL U1812 ( .A0(n3119), .A1(n3256), .B0(n3258), .B1(n819), .Y(n1442) );
  OAI22XL U1813 ( .A0(n3165), .A1(n3255), .B0(n3253), .B1(n810), .Y(n1451) );
  OAI22XL U1814 ( .A0(n3163), .A1(n3255), .B0(n3253), .B1(n809), .Y(n1452) );
  OAI22XL U1815 ( .A0(n3161), .A1(n3255), .B0(n3253), .B1(n808), .Y(n1453) );
  OAI22XL U1816 ( .A0(n3159), .A1(n3255), .B0(n3253), .B1(n807), .Y(n1454) );
  OAI22XL U1817 ( .A0(n3157), .A1(n3252), .B0(n3253), .B1(n806), .Y(n1455) );
  OAI22XL U1818 ( .A0(n3155), .A1(n3255), .B0(n3253), .B1(n805), .Y(n1456) );
  OAI22XL U1819 ( .A0(n3153), .A1(n3252), .B0(n3253), .B1(n804), .Y(n1457) );
  OAI22XL U1820 ( .A0(n3151), .A1(n3252), .B0(n3253), .B1(n803), .Y(n1458) );
  OAI22XL U1821 ( .A0(n3149), .A1(n3255), .B0(n3253), .B1(n802), .Y(n1459) );
  OAI22XL U1822 ( .A0(n3147), .A1(n3255), .B0(n3253), .B1(n801), .Y(n1460) );
  OAI22XL U1823 ( .A0(n3145), .A1(n3252), .B0(n3253), .B1(n800), .Y(n1461) );
  OAI22XL U1824 ( .A0(n3143), .A1(n3255), .B0(n3253), .B1(n799), .Y(n1462) );
  OAI22XL U1825 ( .A0(n3141), .A1(n3252), .B0(n3254), .B1(n798), .Y(n1463) );
  OAI22XL U1826 ( .A0(n3139), .A1(n3252), .B0(n3254), .B1(n797), .Y(n1464) );
  OAI22XL U1827 ( .A0(n3137), .A1(n3252), .B0(n3254), .B1(n796), .Y(n1465) );
  OAI22XL U1828 ( .A0(n3135), .A1(n3252), .B0(n3254), .B1(n795), .Y(n1466) );
  OAI22XL U1829 ( .A0(n3133), .A1(n72), .B0(n3254), .B1(n794), .Y(n1467) );
  OAI22XL U1830 ( .A0(n3131), .A1(n72), .B0(n3254), .B1(n793), .Y(n1468) );
  OAI22XL U1831 ( .A0(n3129), .A1(n72), .B0(n3254), .B1(n792), .Y(n1469) );
  OAI22XL U1832 ( .A0(n3127), .A1(n72), .B0(n3254), .B1(n791), .Y(n1470) );
  OAI22XL U1833 ( .A0(n3125), .A1(n72), .B0(n3254), .B1(n790), .Y(n1471) );
  OAI22XL U1834 ( .A0(n3123), .A1(n3252), .B0(n3254), .B1(n789), .Y(n1472) );
  OAI22XL U1835 ( .A0(n3121), .A1(n3252), .B0(n3254), .B1(n788), .Y(n1473) );
  OAI22XL U1836 ( .A0(n3119), .A1(n3252), .B0(n3254), .B1(n787), .Y(n1474) );
  OAI22XL U1837 ( .A0(n3165), .A1(n3251), .B0(n3249), .B1(n778), .Y(n1483) );
  OAI22XL U1838 ( .A0(n3163), .A1(n3251), .B0(n3249), .B1(n777), .Y(n1484) );
  OAI22XL U1839 ( .A0(n3161), .A1(n3251), .B0(n3249), .B1(n776), .Y(n1485) );
  OAI22XL U1840 ( .A0(n3159), .A1(n3251), .B0(n3249), .B1(n775), .Y(n1486) );
  OAI22XL U1841 ( .A0(n3157), .A1(n3248), .B0(n3249), .B1(n774), .Y(n1487) );
  OAI22XL U1842 ( .A0(n3155), .A1(n3251), .B0(n3249), .B1(n773), .Y(n1488) );
  OAI22XL U1843 ( .A0(n3153), .A1(n3248), .B0(n3249), .B1(n772), .Y(n1489) );
  OAI22XL U1844 ( .A0(n3151), .A1(n3248), .B0(n3249), .B1(n771), .Y(n1490) );
  OAI22XL U1845 ( .A0(n3149), .A1(n3251), .B0(n3249), .B1(n770), .Y(n1491) );
  OAI22XL U1846 ( .A0(n3147), .A1(n3251), .B0(n3249), .B1(n769), .Y(n1492) );
  OAI22XL U1847 ( .A0(n3145), .A1(n3248), .B0(n3249), .B1(n768), .Y(n1493) );
  OAI22XL U1848 ( .A0(n3143), .A1(n3251), .B0(n3249), .B1(n767), .Y(n1494) );
  OAI22XL U1849 ( .A0(n3141), .A1(n3248), .B0(n3250), .B1(n766), .Y(n1495) );
  OAI22XL U1850 ( .A0(n3139), .A1(n3248), .B0(n3250), .B1(n765), .Y(n1496) );
  OAI22XL U1851 ( .A0(n3137), .A1(n3248), .B0(n3250), .B1(n764), .Y(n1497) );
  OAI22XL U1852 ( .A0(n3135), .A1(n3248), .B0(n3250), .B1(n763), .Y(n1498) );
  OAI22XL U1853 ( .A0(n3133), .A1(n74), .B0(n3250), .B1(n762), .Y(n1499) );
  OAI22XL U1854 ( .A0(n3131), .A1(n74), .B0(n3250), .B1(n761), .Y(n1500) );
  OAI22XL U1855 ( .A0(n3129), .A1(n74), .B0(n3250), .B1(n760), .Y(n1501) );
  OAI22XL U1856 ( .A0(n3127), .A1(n74), .B0(n3250), .B1(n759), .Y(n1502) );
  OAI22XL U1857 ( .A0(n3125), .A1(n74), .B0(n3250), .B1(n758), .Y(n1503) );
  OAI22XL U1858 ( .A0(n3123), .A1(n3248), .B0(n3250), .B1(n757), .Y(n1504) );
  OAI22XL U1859 ( .A0(n3121), .A1(n3248), .B0(n3250), .B1(n756), .Y(n1505) );
  OAI22XL U1860 ( .A0(n3119), .A1(n3248), .B0(n3250), .B1(n755), .Y(n1506) );
  OAI22XL U1861 ( .A0(n3165), .A1(n3247), .B0(n3245), .B1(n746), .Y(n1515) );
  OAI22XL U1862 ( .A0(n3163), .A1(n3247), .B0(n3245), .B1(n745), .Y(n1516) );
  OAI22XL U1863 ( .A0(n3161), .A1(n3247), .B0(n3245), .B1(n744), .Y(n1517) );
  OAI22XL U1864 ( .A0(n3159), .A1(n3247), .B0(n3245), .B1(n743), .Y(n1518) );
  OAI22XL U1865 ( .A0(n3157), .A1(n3244), .B0(n3245), .B1(n742), .Y(n1519) );
  OAI22XL U1866 ( .A0(n3155), .A1(n3247), .B0(n3245), .B1(n741), .Y(n1520) );
  OAI22XL U1867 ( .A0(n3153), .A1(n3244), .B0(n3245), .B1(n740), .Y(n1521) );
  OAI22XL U1868 ( .A0(n3151), .A1(n3244), .B0(n3245), .B1(n739), .Y(n1522) );
  OAI22XL U1869 ( .A0(n3149), .A1(n3247), .B0(n3245), .B1(n738), .Y(n1523) );
  OAI22XL U1870 ( .A0(n3147), .A1(n3247), .B0(n3245), .B1(n737), .Y(n1524) );
  OAI22XL U1871 ( .A0(n3145), .A1(n3244), .B0(n3245), .B1(n736), .Y(n1525) );
  OAI22XL U1872 ( .A0(n3143), .A1(n3247), .B0(n3245), .B1(n735), .Y(n1526) );
  OAI22XL U1873 ( .A0(n3141), .A1(n3244), .B0(n3246), .B1(n734), .Y(n1527) );
  OAI22XL U1874 ( .A0(n3139), .A1(n3244), .B0(n3246), .B1(n733), .Y(n1528) );
  OAI22XL U1875 ( .A0(n3137), .A1(n3244), .B0(n3246), .B1(n732), .Y(n1529) );
  OAI22XL U1876 ( .A0(n3135), .A1(n3244), .B0(n3246), .B1(n731), .Y(n1530) );
  OAI22XL U1877 ( .A0(n3133), .A1(n76), .B0(n3246), .B1(n730), .Y(n1531) );
  OAI22XL U1878 ( .A0(n3131), .A1(n76), .B0(n3246), .B1(n729), .Y(n1532) );
  OAI22XL U1879 ( .A0(n3129), .A1(n76), .B0(n3246), .B1(n728), .Y(n1533) );
  OAI22XL U1880 ( .A0(n3127), .A1(n76), .B0(n3246), .B1(n727), .Y(n1534) );
  OAI22XL U1881 ( .A0(n3125), .A1(n76), .B0(n3246), .B1(n726), .Y(n1535) );
  OAI22XL U1882 ( .A0(n3123), .A1(n3244), .B0(n3246), .B1(n725), .Y(n1536) );
  OAI22XL U1883 ( .A0(n3121), .A1(n3244), .B0(n3246), .B1(n724), .Y(n1537) );
  OAI22XL U1884 ( .A0(n3119), .A1(n3244), .B0(n3246), .B1(n723), .Y(n1538) );
  OAI22XL U1885 ( .A0(n3165), .A1(n3243), .B0(n3241), .B1(n714), .Y(n1547) );
  OAI22XL U1886 ( .A0(n3163), .A1(n3243), .B0(n3241), .B1(n713), .Y(n1548) );
  OAI22XL U1887 ( .A0(n3161), .A1(n3243), .B0(n3241), .B1(n712), .Y(n1549) );
  OAI22XL U1888 ( .A0(n3159), .A1(n3243), .B0(n3241), .B1(n711), .Y(n1550) );
  OAI22XL U1889 ( .A0(n3157), .A1(n3240), .B0(n3241), .B1(n710), .Y(n1551) );
  OAI22XL U1890 ( .A0(n3155), .A1(n3243), .B0(n3241), .B1(n709), .Y(n1552) );
  OAI22XL U1891 ( .A0(n3153), .A1(n3240), .B0(n3241), .B1(n708), .Y(n1553) );
  OAI22XL U1892 ( .A0(n3151), .A1(n3240), .B0(n3241), .B1(n707), .Y(n1554) );
  OAI22XL U1893 ( .A0(n3149), .A1(n3243), .B0(n3241), .B1(n706), .Y(n1555) );
  OAI22XL U1894 ( .A0(n3147), .A1(n3243), .B0(n3241), .B1(n705), .Y(n1556) );
  OAI22XL U1895 ( .A0(n3145), .A1(n3240), .B0(n3241), .B1(n704), .Y(n1557) );
  OAI22XL U1896 ( .A0(n3143), .A1(n3243), .B0(n3241), .B1(n703), .Y(n1558) );
  OAI22XL U1897 ( .A0(n3141), .A1(n3240), .B0(n3242), .B1(n702), .Y(n1559) );
  OAI22XL U1898 ( .A0(n3139), .A1(n3240), .B0(n3242), .B1(n701), .Y(n1560) );
  OAI22XL U1899 ( .A0(n3137), .A1(n3240), .B0(n3242), .B1(n700), .Y(n1561) );
  OAI22XL U1900 ( .A0(n3135), .A1(n3240), .B0(n3242), .B1(n699), .Y(n1562) );
  OAI22XL U1901 ( .A0(n3133), .A1(n78), .B0(n3242), .B1(n698), .Y(n1563) );
  OAI22XL U1902 ( .A0(n3131), .A1(n78), .B0(n3242), .B1(n697), .Y(n1564) );
  OAI22XL U1903 ( .A0(n3129), .A1(n78), .B0(n3242), .B1(n696), .Y(n1565) );
  OAI22XL U1904 ( .A0(n3127), .A1(n78), .B0(n3242), .B1(n695), .Y(n1566) );
  OAI22XL U1905 ( .A0(n3125), .A1(n78), .B0(n3242), .B1(n694), .Y(n1567) );
  OAI22XL U1906 ( .A0(n3123), .A1(n3240), .B0(n3242), .B1(n693), .Y(n1568) );
  OAI22XL U1907 ( .A0(n3121), .A1(n3240), .B0(n3242), .B1(n692), .Y(n1569) );
  OAI22XL U1908 ( .A0(n3119), .A1(n3240), .B0(n3242), .B1(n691), .Y(n1570) );
  OAI22XL U1909 ( .A0(n3165), .A1(n3239), .B0(n3237), .B1(n682), .Y(n1579) );
  OAI22XL U1910 ( .A0(n3163), .A1(n3239), .B0(n3237), .B1(n681), .Y(n1580) );
  OAI22XL U1911 ( .A0(n3161), .A1(n3239), .B0(n3237), .B1(n680), .Y(n1581) );
  OAI22XL U1912 ( .A0(n3159), .A1(n3239), .B0(n3237), .B1(n679), .Y(n1582) );
  OAI22XL U1913 ( .A0(n3157), .A1(n3236), .B0(n3237), .B1(n678), .Y(n1583) );
  OAI22XL U1914 ( .A0(n3155), .A1(n3239), .B0(n3237), .B1(n677), .Y(n1584) );
  OAI22XL U1915 ( .A0(n3153), .A1(n3236), .B0(n3237), .B1(n676), .Y(n1585) );
  OAI22XL U1916 ( .A0(n3151), .A1(n3236), .B0(n3237), .B1(n675), .Y(n1586) );
  OAI22XL U1917 ( .A0(n3149), .A1(n3239), .B0(n3237), .B1(n674), .Y(n1587) );
  OAI22XL U1918 ( .A0(n3147), .A1(n3239), .B0(n3237), .B1(n673), .Y(n1588) );
  OAI22XL U1919 ( .A0(n3145), .A1(n3236), .B0(n3237), .B1(n672), .Y(n1589) );
  OAI22XL U1920 ( .A0(n3143), .A1(n3239), .B0(n3237), .B1(n671), .Y(n1590) );
  OAI22XL U1921 ( .A0(n3141), .A1(n3236), .B0(n3238), .B1(n670), .Y(n1591) );
  OAI22XL U1922 ( .A0(n3139), .A1(n3236), .B0(n3238), .B1(n669), .Y(n1592) );
  OAI22XL U1923 ( .A0(n3137), .A1(n3236), .B0(n3238), .B1(n668), .Y(n1593) );
  OAI22XL U1924 ( .A0(n3135), .A1(n3236), .B0(n3238), .B1(n667), .Y(n1594) );
  OAI22XL U1925 ( .A0(n3133), .A1(n81), .B0(n3238), .B1(n666), .Y(n1595) );
  OAI22XL U1926 ( .A0(n3131), .A1(n81), .B0(n3238), .B1(n665), .Y(n1596) );
  OAI22XL U1927 ( .A0(n3129), .A1(n81), .B0(n3238), .B1(n664), .Y(n1597) );
  OAI22XL U1928 ( .A0(n3127), .A1(n81), .B0(n3238), .B1(n663), .Y(n1598) );
  OAI22XL U1929 ( .A0(n3125), .A1(n81), .B0(n3238), .B1(n662), .Y(n1599) );
  OAI22XL U1930 ( .A0(n3123), .A1(n3236), .B0(n3238), .B1(n661), .Y(n1600) );
  OAI22XL U1931 ( .A0(n3121), .A1(n3236), .B0(n3238), .B1(n660), .Y(n1601) );
  OAI22XL U1932 ( .A0(n3119), .A1(n3236), .B0(n3238), .B1(n659), .Y(n1602) );
  OAI22XL U1933 ( .A0(n3165), .A1(n3235), .B0(n3233), .B1(n650), .Y(n1611) );
  OAI22XL U1934 ( .A0(n3163), .A1(n3235), .B0(n3233), .B1(n649), .Y(n1612) );
  OAI22XL U1935 ( .A0(n3161), .A1(n3235), .B0(n3233), .B1(n648), .Y(n1613) );
  OAI22XL U1936 ( .A0(n3159), .A1(n3235), .B0(n3233), .B1(n647), .Y(n1614) );
  OAI22XL U1937 ( .A0(n3157), .A1(n3235), .B0(n3233), .B1(n646), .Y(n1615) );
  OAI22XL U1938 ( .A0(n3155), .A1(n3235), .B0(n3233), .B1(n645), .Y(n1616) );
  OAI22XL U1939 ( .A0(n3153), .A1(n3235), .B0(n3233), .B1(n644), .Y(n1617) );
  OAI22XL U1940 ( .A0(n3151), .A1(n3232), .B0(n3233), .B1(n643), .Y(n1618) );
  OAI22XL U1941 ( .A0(n3149), .A1(n3235), .B0(n3233), .B1(n642), .Y(n1619) );
  OAI22XL U1942 ( .A0(n3147), .A1(n3235), .B0(n3233), .B1(n641), .Y(n1620) );
  OAI22XL U1943 ( .A0(n3145), .A1(n3235), .B0(n3233), .B1(n640), .Y(n1621) );
  OAI22XL U1944 ( .A0(n3143), .A1(n3235), .B0(n3233), .B1(n639), .Y(n1622) );
  OAI22XL U1945 ( .A0(n3141), .A1(n3232), .B0(n3234), .B1(n638), .Y(n1623) );
  OAI22XL U1946 ( .A0(n3139), .A1(n3232), .B0(n3234), .B1(n637), .Y(n1624) );
  OAI22XL U1947 ( .A0(n3137), .A1(n3232), .B0(n3234), .B1(n636), .Y(n1625) );
  OAI22XL U1948 ( .A0(n3135), .A1(n3232), .B0(n3234), .B1(n635), .Y(n1626) );
  OAI22XL U1949 ( .A0(n3133), .A1(n3232), .B0(n3234), .B1(n634), .Y(n1627) );
  OAI22XL U1950 ( .A0(n3131), .A1(n3235), .B0(n3234), .B1(n633), .Y(n1628) );
  OAI22XL U1951 ( .A0(n3129), .A1(n3232), .B0(n3234), .B1(n632), .Y(n1629) );
  OAI22XL U1952 ( .A0(n3127), .A1(n3235), .B0(n3234), .B1(n631), .Y(n1630) );
  OAI22XL U1953 ( .A0(n3125), .A1(n3232), .B0(n3234), .B1(n630), .Y(n1631) );
  OAI22XL U1954 ( .A0(n3123), .A1(n3232), .B0(n3234), .B1(n629), .Y(n1632) );
  OAI22XL U1955 ( .A0(n3121), .A1(n3235), .B0(n3234), .B1(n628), .Y(n1633) );
  OAI22XL U1956 ( .A0(n3119), .A1(n3235), .B0(n3234), .B1(n627), .Y(n1634) );
  OAI22XL U1957 ( .A0(n3165), .A1(n3231), .B0(n3229), .B1(n618), .Y(n1643) );
  OAI22XL U1958 ( .A0(n3163), .A1(n3231), .B0(n3229), .B1(n617), .Y(n1644) );
  OAI22XL U1959 ( .A0(n3161), .A1(n3231), .B0(n3229), .B1(n616), .Y(n1645) );
  OAI22XL U1960 ( .A0(n3159), .A1(n3231), .B0(n3229), .B1(n615), .Y(n1646) );
  OAI22XL U1961 ( .A0(n3157), .A1(n3231), .B0(n3229), .B1(n614), .Y(n1647) );
  OAI22XL U1962 ( .A0(n3155), .A1(n3231), .B0(n3229), .B1(n613), .Y(n1648) );
  OAI22XL U1963 ( .A0(n3153), .A1(n3231), .B0(n3229), .B1(n612), .Y(n1649) );
  OAI22XL U1964 ( .A0(n3151), .A1(n3228), .B0(n3229), .B1(n611), .Y(n1650) );
  OAI22XL U1965 ( .A0(n3149), .A1(n3231), .B0(n3229), .B1(n610), .Y(n1651) );
  OAI22XL U1966 ( .A0(n3147), .A1(n3231), .B0(n3229), .B1(n609), .Y(n1652) );
  OAI22XL U1967 ( .A0(n3145), .A1(n3231), .B0(n3229), .B1(n608), .Y(n1653) );
  OAI22XL U1968 ( .A0(n3143), .A1(n3231), .B0(n3229), .B1(n607), .Y(n1654) );
  OAI22XL U1969 ( .A0(n3141), .A1(n3228), .B0(n3230), .B1(n606), .Y(n1655) );
  OAI22XL U1970 ( .A0(n3139), .A1(n3228), .B0(n3230), .B1(n605), .Y(n1656) );
  OAI22XL U1971 ( .A0(n3137), .A1(n3228), .B0(n3230), .B1(n604), .Y(n1657) );
  OAI22XL U1972 ( .A0(n3135), .A1(n3228), .B0(n3230), .B1(n603), .Y(n1658) );
  OAI22XL U1973 ( .A0(n3133), .A1(n3228), .B0(n3230), .B1(n602), .Y(n1659) );
  OAI22XL U1974 ( .A0(n3131), .A1(n3231), .B0(n3230), .B1(n601), .Y(n1660) );
  OAI22XL U1975 ( .A0(n3129), .A1(n3228), .B0(n3230), .B1(n600), .Y(n1661) );
  OAI22XL U1976 ( .A0(n3127), .A1(n3231), .B0(n3230), .B1(n599), .Y(n1662) );
  OAI22XL U1977 ( .A0(n3125), .A1(n3228), .B0(n3230), .B1(n598), .Y(n1663) );
  OAI22XL U1978 ( .A0(n3123), .A1(n3228), .B0(n3230), .B1(n597), .Y(n1664) );
  OAI22XL U1979 ( .A0(n3121), .A1(n3231), .B0(n3230), .B1(n596), .Y(n1665) );
  OAI22XL U1980 ( .A0(n3119), .A1(n3231), .B0(n3230), .B1(n595), .Y(n1666) );
  OAI22XL U1981 ( .A0(n3165), .A1(n3227), .B0(n3225), .B1(n586), .Y(n1675) );
  OAI22XL U1982 ( .A0(n3163), .A1(n3227), .B0(n3225), .B1(n585), .Y(n1676) );
  OAI22XL U1983 ( .A0(n3161), .A1(n3227), .B0(n3225), .B1(n584), .Y(n1677) );
  OAI22XL U1984 ( .A0(n3159), .A1(n3227), .B0(n3225), .B1(n583), .Y(n1678) );
  OAI22XL U1985 ( .A0(n3157), .A1(n3227), .B0(n3225), .B1(n582), .Y(n1679) );
  OAI22XL U1986 ( .A0(n3155), .A1(n3227), .B0(n3225), .B1(n581), .Y(n1680) );
  OAI22XL U1987 ( .A0(n3153), .A1(n3227), .B0(n3225), .B1(n580), .Y(n1681) );
  OAI22XL U1988 ( .A0(n3151), .A1(n3224), .B0(n3225), .B1(n579), .Y(n1682) );
  OAI22XL U1989 ( .A0(n3149), .A1(n3227), .B0(n3225), .B1(n578), .Y(n1683) );
  OAI22XL U1990 ( .A0(n3147), .A1(n3227), .B0(n3225), .B1(n577), .Y(n1684) );
  OAI22XL U1991 ( .A0(n3145), .A1(n3227), .B0(n3225), .B1(n576), .Y(n1685) );
  OAI22XL U1992 ( .A0(n3143), .A1(n3227), .B0(n3225), .B1(n575), .Y(n1686) );
  OAI22XL U1993 ( .A0(n3141), .A1(n3224), .B0(n3226), .B1(n574), .Y(n1687) );
  OAI22XL U1994 ( .A0(n3139), .A1(n3224), .B0(n3226), .B1(n573), .Y(n1688) );
  OAI22XL U1995 ( .A0(n3137), .A1(n3224), .B0(n3226), .B1(n572), .Y(n1689) );
  OAI22XL U1996 ( .A0(n3135), .A1(n3224), .B0(n3226), .B1(n571), .Y(n1690) );
  OAI22XL U1997 ( .A0(n3133), .A1(n3224), .B0(n3226), .B1(n570), .Y(n1691) );
  OAI22XL U1998 ( .A0(n3131), .A1(n3227), .B0(n3226), .B1(n569), .Y(n1692) );
  OAI22XL U1999 ( .A0(n3129), .A1(n3224), .B0(n3226), .B1(n568), .Y(n1693) );
  OAI22XL U2000 ( .A0(n3127), .A1(n3227), .B0(n3226), .B1(n567), .Y(n1694) );
  OAI22XL U2001 ( .A0(n3125), .A1(n3224), .B0(n3226), .B1(n566), .Y(n1695) );
  OAI22XL U2002 ( .A0(n3123), .A1(n3224), .B0(n3226), .B1(n565), .Y(n1696) );
  OAI22XL U2003 ( .A0(n3121), .A1(n3227), .B0(n3226), .B1(n564), .Y(n1697) );
  OAI22XL U2004 ( .A0(n3119), .A1(n3227), .B0(n3226), .B1(n563), .Y(n1698) );
  OAI22XL U2005 ( .A0(n3165), .A1(n3223), .B0(n3221), .B1(n554), .Y(n1707) );
  OAI22XL U2006 ( .A0(n3163), .A1(n3223), .B0(n3221), .B1(n553), .Y(n1708) );
  OAI22XL U2007 ( .A0(n3161), .A1(n3223), .B0(n3221), .B1(n552), .Y(n1709) );
  OAI22XL U2008 ( .A0(n3159), .A1(n3223), .B0(n3221), .B1(n551), .Y(n1710) );
  OAI22XL U2009 ( .A0(n3157), .A1(n3223), .B0(n3221), .B1(n550), .Y(n1711) );
  OAI22XL U2010 ( .A0(n3155), .A1(n3223), .B0(n3221), .B1(n549), .Y(n1712) );
  OAI22XL U2011 ( .A0(n3153), .A1(n3223), .B0(n3221), .B1(n548), .Y(n1713) );
  OAI22XL U2012 ( .A0(n3151), .A1(n3220), .B0(n3221), .B1(n547), .Y(n1714) );
  OAI22XL U2013 ( .A0(n3149), .A1(n3223), .B0(n3221), .B1(n546), .Y(n1715) );
  OAI22XL U2014 ( .A0(n3147), .A1(n3223), .B0(n3221), .B1(n545), .Y(n1716) );
  OAI22XL U2015 ( .A0(n3145), .A1(n3223), .B0(n3221), .B1(n544), .Y(n1717) );
  OAI22XL U2016 ( .A0(n3143), .A1(n3223), .B0(n3221), .B1(n543), .Y(n1718) );
  OAI22XL U2017 ( .A0(n3141), .A1(n3220), .B0(n3222), .B1(n542), .Y(n1719) );
  OAI22XL U2018 ( .A0(n3139), .A1(n3220), .B0(n3222), .B1(n541), .Y(n1720) );
  OAI22XL U2019 ( .A0(n3137), .A1(n3220), .B0(n3222), .B1(n540), .Y(n1721) );
  OAI22XL U2020 ( .A0(n3135), .A1(n3220), .B0(n3222), .B1(n539), .Y(n1722) );
  OAI22XL U2021 ( .A0(n3133), .A1(n3220), .B0(n3222), .B1(n538), .Y(n1723) );
  OAI22XL U2022 ( .A0(n3131), .A1(n3223), .B0(n3222), .B1(n537), .Y(n1724) );
  OAI22XL U2023 ( .A0(n3129), .A1(n3220), .B0(n3222), .B1(n536), .Y(n1725) );
  OAI22XL U2024 ( .A0(n3127), .A1(n3223), .B0(n3222), .B1(n535), .Y(n1726) );
  OAI22XL U2025 ( .A0(n3125), .A1(n3220), .B0(n3222), .B1(n534), .Y(n1727) );
  OAI22XL U2026 ( .A0(n3123), .A1(n3220), .B0(n3222), .B1(n533), .Y(n1728) );
  OAI22XL U2027 ( .A0(n3121), .A1(n3223), .B0(n3222), .B1(n532), .Y(n1729) );
  OAI22XL U2028 ( .A0(n3119), .A1(n3223), .B0(n3222), .B1(n531), .Y(n1730) );
  OAI22XL U2029 ( .A0(n3165), .A1(n3219), .B0(n3217), .B1(n522), .Y(n1739) );
  OAI22XL U2030 ( .A0(n3163), .A1(n3219), .B0(n3217), .B1(n521), .Y(n1740) );
  OAI22XL U2031 ( .A0(n3161), .A1(n3219), .B0(n3217), .B1(n520), .Y(n1741) );
  OAI22XL U2032 ( .A0(n3159), .A1(n3219), .B0(n3217), .B1(n519), .Y(n1742) );
  OAI22XL U2033 ( .A0(n3157), .A1(n3216), .B0(n3217), .B1(n518), .Y(n1743) );
  OAI22XL U2034 ( .A0(n3155), .A1(n3216), .B0(n3217), .B1(n517), .Y(n1744) );
  OAI22XL U2035 ( .A0(n3153), .A1(n3216), .B0(n3217), .B1(n516), .Y(n1745) );
  OAI22XL U2036 ( .A0(n3151), .A1(n3216), .B0(n3217), .B1(n515), .Y(n1746) );
  OAI22XL U2037 ( .A0(n3149), .A1(n3216), .B0(n3217), .B1(n514), .Y(n1747) );
  OAI22XL U2038 ( .A0(n3147), .A1(n3216), .B0(n3217), .B1(n513), .Y(n1748) );
  OAI22XL U2039 ( .A0(n3145), .A1(n3216), .B0(n3217), .B1(n512), .Y(n1749) );
  OAI22XL U2040 ( .A0(n3143), .A1(n3219), .B0(n3217), .B1(n511), .Y(n1750) );
  OAI22XL U2041 ( .A0(n3141), .A1(n3216), .B0(n3218), .B1(n510), .Y(n1751) );
  OAI22XL U2042 ( .A0(n3139), .A1(n3216), .B0(n3218), .B1(n509), .Y(n1752) );
  OAI22XL U2043 ( .A0(n3137), .A1(n94), .B0(n3218), .B1(n508), .Y(n1753) );
  OAI22XL U2044 ( .A0(n3135), .A1(n3216), .B0(n3217), .B1(n507), .Y(n1754) );
  OAI22XL U2045 ( .A0(n3133), .A1(n3219), .B0(n3218), .B1(n506), .Y(n1755) );
  OAI22XL U2046 ( .A0(n3131), .A1(n3219), .B0(n3217), .B1(n505), .Y(n1756) );
  OAI22XL U2047 ( .A0(n3129), .A1(n3216), .B0(n3218), .B1(n504), .Y(n1757) );
  OAI22XL U2048 ( .A0(n3127), .A1(n3219), .B0(n3217), .B1(n503), .Y(n1758) );
  OAI22XL U2049 ( .A0(n3125), .A1(n3216), .B0(n3218), .B1(n502), .Y(n1759) );
  OAI22XL U2050 ( .A0(n3123), .A1(n3216), .B0(n3217), .B1(n501), .Y(n1760) );
  OAI22XL U2051 ( .A0(n3121), .A1(n94), .B0(n3218), .B1(n500), .Y(n1761) );
  OAI22XL U2052 ( .A0(n3119), .A1(n3219), .B0(n3217), .B1(n499), .Y(n1762) );
  OAI22XL U2053 ( .A0(n3164), .A1(n3212), .B0(n3214), .B1(n490), .Y(n1771) );
  OAI22XL U2054 ( .A0(n3162), .A1(n3212), .B0(n3214), .B1(n489), .Y(n1772) );
  OAI22XL U2055 ( .A0(n3160), .A1(n3212), .B0(n3214), .B1(n488), .Y(n1773) );
  OAI22XL U2056 ( .A0(n3158), .A1(n3212), .B0(n3214), .B1(n487), .Y(n1774) );
  OAI22XL U2057 ( .A0(n3156), .A1(n3212), .B0(n3214), .B1(n486), .Y(n1775) );
  OAI22XL U2058 ( .A0(n3154), .A1(n3212), .B0(n3214), .B1(n485), .Y(n1776) );
  OAI22XL U2059 ( .A0(n3152), .A1(n3212), .B0(n3214), .B1(n484), .Y(n1777) );
  OAI22XL U2060 ( .A0(n3150), .A1(n3213), .B0(n3214), .B1(n483), .Y(n1778) );
  OAI22XL U2061 ( .A0(n3148), .A1(n3212), .B0(n3214), .B1(n482), .Y(n1779) );
  OAI22XL U2062 ( .A0(n3146), .A1(n3212), .B0(n3214), .B1(n481), .Y(n1780) );
  OAI22XL U2063 ( .A0(n3144), .A1(n3212), .B0(n3214), .B1(n480), .Y(n1781) );
  OAI22XL U2064 ( .A0(n3142), .A1(n3213), .B0(n3214), .B1(n479), .Y(n1782) );
  OAI22XL U2065 ( .A0(n3140), .A1(n3213), .B0(n3215), .B1(n478), .Y(n1783) );
  OAI22XL U2066 ( .A0(n3138), .A1(n3213), .B0(n3215), .B1(n477), .Y(n1784) );
  OAI22XL U2067 ( .A0(n3136), .A1(n3213), .B0(n3215), .B1(n476), .Y(n1785) );
  OAI22XL U2068 ( .A0(n3134), .A1(n3213), .B0(n3215), .B1(n475), .Y(n1786) );
  OAI22XL U2069 ( .A0(n3132), .A1(n3213), .B0(n3215), .B1(n474), .Y(n1787) );
  OAI22XL U2070 ( .A0(n3130), .A1(n96), .B0(n3215), .B1(n473), .Y(n1788) );
  OAI22XL U2071 ( .A0(n3128), .A1(n3213), .B0(n3215), .B1(n472), .Y(n1789) );
  OAI22XL U2072 ( .A0(n3126), .A1(n96), .B0(n3215), .B1(n471), .Y(n1790) );
  OAI22XL U2073 ( .A0(n3124), .A1(n3213), .B0(n3215), .B1(n470), .Y(n1791) );
  OAI22XL U2074 ( .A0(n3122), .A1(n3212), .B0(n3215), .B1(n469), .Y(n1792) );
  OAI22XL U2075 ( .A0(n3120), .A1(n3213), .B0(n3215), .B1(n468), .Y(n1793) );
  OAI22XL U2076 ( .A0(n3118), .A1(n3213), .B0(n3215), .B1(n467), .Y(n1794) );
  OAI22XL U2077 ( .A0(n3164), .A1(n3208), .B0(n3210), .B1(n458), .Y(n1803) );
  OAI22XL U2078 ( .A0(n3162), .A1(n3208), .B0(n3210), .B1(n457), .Y(n1804) );
  OAI22XL U2079 ( .A0(n3160), .A1(n3208), .B0(n3210), .B1(n456), .Y(n1805) );
  OAI22XL U2080 ( .A0(n3158), .A1(n3208), .B0(n3210), .B1(n455), .Y(n1806) );
  OAI22XL U2081 ( .A0(n3156), .A1(n3208), .B0(n3210), .B1(n454), .Y(n1807) );
  OAI22XL U2082 ( .A0(n3154), .A1(n3208), .B0(n3210), .B1(n453), .Y(n1808) );
  OAI22XL U2083 ( .A0(n3152), .A1(n3208), .B0(n3210), .B1(n452), .Y(n1809) );
  OAI22XL U2084 ( .A0(n3150), .A1(n3209), .B0(n3210), .B1(n451), .Y(n1810) );
  OAI22XL U2085 ( .A0(n3148), .A1(n3208), .B0(n3210), .B1(n450), .Y(n1811) );
  OAI22XL U2086 ( .A0(n3146), .A1(n3208), .B0(n3210), .B1(n449), .Y(n1812) );
  OAI22XL U2087 ( .A0(n3144), .A1(n3208), .B0(n3210), .B1(n448), .Y(n1813) );
  OAI22XL U2088 ( .A0(n3142), .A1(n3209), .B0(n3210), .B1(n447), .Y(n1814) );
  OAI22XL U2089 ( .A0(n3140), .A1(n3209), .B0(n3211), .B1(n446), .Y(n1815) );
  OAI22XL U2090 ( .A0(n3138), .A1(n3209), .B0(n3211), .B1(n445), .Y(n1816) );
  OAI22XL U2091 ( .A0(n3136), .A1(n3209), .B0(n3211), .B1(n444), .Y(n1817) );
  OAI22XL U2092 ( .A0(n3134), .A1(n3209), .B0(n3211), .B1(n443), .Y(n1818) );
  OAI22XL U2093 ( .A0(n3132), .A1(n3209), .B0(n3211), .B1(n442), .Y(n1819) );
  OAI22XL U2094 ( .A0(n3130), .A1(n98), .B0(n3211), .B1(n441), .Y(n1820) );
  OAI22XL U2095 ( .A0(n3128), .A1(n3209), .B0(n3211), .B1(n440), .Y(n1821) );
  OAI22XL U2096 ( .A0(n3126), .A1(n98), .B0(n3211), .B1(n439), .Y(n1822) );
  OAI22XL U2097 ( .A0(n3124), .A1(n3209), .B0(n3211), .B1(n438), .Y(n1823) );
  OAI22XL U2098 ( .A0(n3122), .A1(n3208), .B0(n3211), .B1(n437), .Y(n1824) );
  OAI22XL U2099 ( .A0(n3120), .A1(n3209), .B0(n3211), .B1(n436), .Y(n1825) );
  OAI22XL U2100 ( .A0(n3118), .A1(n3209), .B0(n3211), .B1(n435), .Y(n1826) );
  OAI22XL U2101 ( .A0(n3164), .A1(n3207), .B0(n3205), .B1(n426), .Y(n1835) );
  OAI22XL U2102 ( .A0(n3162), .A1(n3207), .B0(n3205), .B1(n425), .Y(n1836) );
  OAI22XL U2103 ( .A0(n3160), .A1(n3207), .B0(n3205), .B1(n424), .Y(n1837) );
  OAI22XL U2104 ( .A0(n3158), .A1(n3207), .B0(n3205), .B1(n423), .Y(n1838) );
  OAI22XL U2105 ( .A0(n3156), .A1(n3204), .B0(n3205), .B1(n422), .Y(n1839) );
  OAI22XL U2106 ( .A0(n3154), .A1(n101), .B0(n3205), .B1(n421), .Y(n1840) );
  OAI22XL U2107 ( .A0(n3152), .A1(n101), .B0(n3205), .B1(n420), .Y(n1841) );
  OAI22XL U2108 ( .A0(n3150), .A1(n3207), .B0(n3205), .B1(n419), .Y(n1842) );
  OAI22XL U2109 ( .A0(n3148), .A1(n3207), .B0(n3205), .B1(n418), .Y(n1843) );
  OAI22XL U2110 ( .A0(n3146), .A1(n3207), .B0(n3205), .B1(n417), .Y(n1844) );
  OAI22XL U2111 ( .A0(n3144), .A1(n3207), .B0(n3205), .B1(n416), .Y(n1845) );
  OAI22XL U2112 ( .A0(n3142), .A1(n3204), .B0(n3205), .B1(n415), .Y(n1846) );
  OAI22XL U2113 ( .A0(n3140), .A1(n3204), .B0(n3206), .B1(n414), .Y(n1847) );
  OAI22XL U2114 ( .A0(n3138), .A1(n3204), .B0(n3205), .B1(n413), .Y(n1848) );
  OAI22XL U2115 ( .A0(n3136), .A1(n3204), .B0(n3206), .B1(n412), .Y(n1849) );
  OAI22XL U2116 ( .A0(n3134), .A1(n3204), .B0(n3205), .B1(n411), .Y(n1850) );
  OAI22XL U2117 ( .A0(n3132), .A1(n3207), .B0(n3206), .B1(n410), .Y(n1851) );
  OAI22XL U2118 ( .A0(n3130), .A1(n3204), .B0(n3205), .B1(n409), .Y(n1852) );
  OAI22XL U2119 ( .A0(n3128), .A1(n3204), .B0(n3206), .B1(n408), .Y(n1853) );
  OAI22XL U2120 ( .A0(n3126), .A1(n3207), .B0(n3205), .B1(n407), .Y(n1854) );
  OAI22XL U2121 ( .A0(n3124), .A1(n3204), .B0(n3206), .B1(n406), .Y(n1855) );
  OAI22XL U2122 ( .A0(n3122), .A1(n3204), .B0(n3205), .B1(n405), .Y(n1856) );
  OAI22XL U2123 ( .A0(n3120), .A1(n3207), .B0(n3206), .B1(n404), .Y(n1857) );
  OAI22XL U2124 ( .A0(n3118), .A1(n3207), .B0(n3205), .B1(n403), .Y(n1858) );
  OAI22XL U2125 ( .A0(n3164), .A1(n3203), .B0(n3201), .B1(n394), .Y(n1867) );
  OAI22XL U2126 ( .A0(n3162), .A1(n3203), .B0(n3201), .B1(n393), .Y(n1868) );
  OAI22XL U2127 ( .A0(n3160), .A1(n3203), .B0(n3201), .B1(n392), .Y(n1869) );
  OAI22XL U2128 ( .A0(n3158), .A1(n3203), .B0(n3201), .B1(n391), .Y(n1870) );
  OAI22XL U2129 ( .A0(n3156), .A1(n3200), .B0(n3201), .B1(n390), .Y(n1871) );
  OAI22XL U2130 ( .A0(n3154), .A1(n3203), .B0(n3201), .B1(n389), .Y(n1872) );
  OAI22XL U2131 ( .A0(n3152), .A1(n3200), .B0(n3201), .B1(n388), .Y(n1873) );
  OAI22XL U2132 ( .A0(n3150), .A1(n3200), .B0(n3201), .B1(n387), .Y(n1874) );
  OAI22XL U2133 ( .A0(n3148), .A1(n3203), .B0(n3201), .B1(n386), .Y(n1875) );
  OAI22XL U2134 ( .A0(n3146), .A1(n3203), .B0(n3201), .B1(n385), .Y(n1876) );
  OAI22XL U2135 ( .A0(n3144), .A1(n3200), .B0(n3201), .B1(n384), .Y(n1877) );
  OAI22XL U2136 ( .A0(n3142), .A1(n3203), .B0(n3201), .B1(n383), .Y(n1878) );
  OAI22XL U2137 ( .A0(n3140), .A1(n3200), .B0(n3202), .B1(n382), .Y(n1879) );
  OAI22XL U2138 ( .A0(n3138), .A1(n3200), .B0(n3202), .B1(n381), .Y(n1880) );
  OAI22XL U2139 ( .A0(n3136), .A1(n3200), .B0(n3202), .B1(n380), .Y(n1881) );
  OAI22XL U2140 ( .A0(n3134), .A1(n3200), .B0(n3202), .B1(n379), .Y(n1882) );
  OAI22XL U2141 ( .A0(n3132), .A1(n104), .B0(n3202), .B1(n378), .Y(n1883) );
  OAI22XL U2142 ( .A0(n3130), .A1(n104), .B0(n3202), .B1(n377), .Y(n1884) );
  OAI22XL U2143 ( .A0(n3128), .A1(n104), .B0(n3202), .B1(n376), .Y(n1885) );
  OAI22XL U2144 ( .A0(n3126), .A1(n104), .B0(n3202), .B1(n375), .Y(n1886) );
  OAI22XL U2145 ( .A0(n3124), .A1(n104), .B0(n3202), .B1(n374), .Y(n1887) );
  OAI22XL U2146 ( .A0(n3122), .A1(n3200), .B0(n3202), .B1(n373), .Y(n1888) );
  OAI22XL U2147 ( .A0(n3120), .A1(n3200), .B0(n3202), .B1(n372), .Y(n1889) );
  OAI22XL U2148 ( .A0(n3118), .A1(n3200), .B0(n3202), .B1(n371), .Y(n1890) );
  OAI22XL U2149 ( .A0(n3164), .A1(n3199), .B0(n3197), .B1(n362), .Y(n1899) );
  OAI22XL U2150 ( .A0(n3162), .A1(n3199), .B0(n3197), .B1(n361), .Y(n1900) );
  OAI22XL U2151 ( .A0(n3160), .A1(n3199), .B0(n3197), .B1(n360), .Y(n1901) );
  OAI22XL U2152 ( .A0(n3158), .A1(n3199), .B0(n3197), .B1(n359), .Y(n1902) );
  OAI22XL U2153 ( .A0(n3156), .A1(n3196), .B0(n3197), .B1(n358), .Y(n1903) );
  OAI22XL U2154 ( .A0(n3154), .A1(n3196), .B0(n3197), .B1(n357), .Y(n1904) );
  OAI22XL U2155 ( .A0(n3152), .A1(n3196), .B0(n3197), .B1(n356), .Y(n1905) );
  OAI22XL U2156 ( .A0(n3150), .A1(n3196), .B0(n3197), .B1(n355), .Y(n1906) );
  OAI22XL U2157 ( .A0(n3148), .A1(n3196), .B0(n3197), .B1(n354), .Y(n1907) );
  OAI22XL U2158 ( .A0(n3146), .A1(n3196), .B0(n3197), .B1(n353), .Y(n1908) );
  OAI22XL U2159 ( .A0(n3144), .A1(n3199), .B0(n3197), .B1(n352), .Y(n1909) );
  OAI22XL U2160 ( .A0(n3142), .A1(n3199), .B0(n3197), .B1(n351), .Y(n1910) );
  OAI22XL U2161 ( .A0(n3140), .A1(n107), .B0(n3198), .B1(n350), .Y(n1911) );
  OAI22XL U2162 ( .A0(n3138), .A1(n107), .B0(n3198), .B1(n349), .Y(n1912) );
  OAI22XL U2163 ( .A0(n3136), .A1(n3196), .B0(n3198), .B1(n348), .Y(n1913) );
  OAI22XL U2164 ( .A0(n3134), .A1(n3196), .B0(n3198), .B1(n347), .Y(n1914) );
  OAI22XL U2165 ( .A0(n3132), .A1(n3196), .B0(n3198), .B1(n346), .Y(n1915) );
  OAI22XL U2166 ( .A0(n3130), .A1(n3196), .B0(n3198), .B1(n345), .Y(n1916) );
  OAI22XL U2167 ( .A0(n3128), .A1(n107), .B0(n3198), .B1(n344), .Y(n1917) );
  OAI22XL U2168 ( .A0(n3126), .A1(n107), .B0(n3198), .B1(n343), .Y(n1918) );
  OAI22XL U2169 ( .A0(n3124), .A1(n3196), .B0(n3198), .B1(n342), .Y(n1919) );
  OAI22XL U2170 ( .A0(n3122), .A1(n3196), .B0(n3198), .B1(n341), .Y(n1920) );
  OAI22XL U2171 ( .A0(n3120), .A1(n3196), .B0(n3198), .B1(n340), .Y(n1921) );
  OAI22XL U2172 ( .A0(n3118), .A1(n3196), .B0(n3198), .B1(n339), .Y(n1922) );
  OAI22XL U2173 ( .A0(n3164), .A1(n3195), .B0(n3193), .B1(n330), .Y(n1931) );
  OAI22XL U2174 ( .A0(n3162), .A1(n3195), .B0(n3193), .B1(n329), .Y(n1932) );
  OAI22XL U2175 ( .A0(n3160), .A1(n3195), .B0(n3193), .B1(n328), .Y(n1933) );
  OAI22XL U2176 ( .A0(n3158), .A1(n3195), .B0(n3193), .B1(n327), .Y(n1934) );
  OAI22XL U2177 ( .A0(n3156), .A1(n3192), .B0(n3193), .B1(n326), .Y(n1935) );
  OAI22XL U2178 ( .A0(n3154), .A1(n3195), .B0(n3193), .B1(n325), .Y(n1936) );
  OAI22XL U2179 ( .A0(n3152), .A1(n3192), .B0(n3193), .B1(n324), .Y(n1937) );
  OAI22XL U2180 ( .A0(n3150), .A1(n3192), .B0(n3193), .B1(n323), .Y(n1938) );
  OAI22XL U2181 ( .A0(n3148), .A1(n3195), .B0(n3193), .B1(n322), .Y(n1939) );
  OAI22XL U2182 ( .A0(n3146), .A1(n3195), .B0(n3193), .B1(n321), .Y(n1940) );
  OAI22XL U2183 ( .A0(n3144), .A1(n3192), .B0(n3193), .B1(n320), .Y(n1941) );
  OAI22XL U2184 ( .A0(n3142), .A1(n3195), .B0(n3193), .B1(n319), .Y(n1942) );
  OAI22XL U2185 ( .A0(n3140), .A1(n3192), .B0(n3194), .B1(n318), .Y(n1943) );
  OAI22XL U2186 ( .A0(n3138), .A1(n3192), .B0(n3194), .B1(n317), .Y(n1944) );
  OAI22XL U2187 ( .A0(n3136), .A1(n3192), .B0(n3194), .B1(n316), .Y(n1945) );
  OAI22XL U2188 ( .A0(n3134), .A1(n3192), .B0(n3194), .B1(n315), .Y(n1946) );
  OAI22XL U2189 ( .A0(n3132), .A1(n110), .B0(n3194), .B1(n314), .Y(n1947) );
  OAI22XL U2190 ( .A0(n3130), .A1(n110), .B0(n3194), .B1(n313), .Y(n1948) );
  OAI22XL U2191 ( .A0(n3128), .A1(n110), .B0(n3194), .B1(n312), .Y(n1949) );
  OAI22XL U2192 ( .A0(n3126), .A1(n110), .B0(n3194), .B1(n311), .Y(n1950) );
  OAI22XL U2193 ( .A0(n3124), .A1(n110), .B0(n3194), .B1(n310), .Y(n1951) );
  OAI22XL U2194 ( .A0(n3122), .A1(n3192), .B0(n3194), .B1(n309), .Y(n1952) );
  OAI22XL U2195 ( .A0(n3120), .A1(n3192), .B0(n3194), .B1(n308), .Y(n1953) );
  OAI22XL U2196 ( .A0(n3118), .A1(n3192), .B0(n3194), .B1(n307), .Y(n1954) );
  OAI22XL U2197 ( .A0(n3164), .A1(n3191), .B0(n3189), .B1(n298), .Y(n1963) );
  OAI22XL U2198 ( .A0(n3162), .A1(n3191), .B0(n3189), .B1(n297), .Y(n1964) );
  OAI22XL U2199 ( .A0(n3160), .A1(n3191), .B0(n3189), .B1(n296), .Y(n1965) );
  OAI22XL U2200 ( .A0(n3158), .A1(n3191), .B0(n3189), .B1(n295), .Y(n1966) );
  OAI22XL U2201 ( .A0(n3156), .A1(n3188), .B0(n3189), .B1(n294), .Y(n1967) );
  OAI22XL U2202 ( .A0(n3154), .A1(n3188), .B0(n3189), .B1(n293), .Y(n1968) );
  OAI22XL U2203 ( .A0(n3152), .A1(n3188), .B0(n3189), .B1(n292), .Y(n1969) );
  OAI22XL U2204 ( .A0(n3150), .A1(n3188), .B0(n3189), .B1(n291), .Y(n1970) );
  OAI22XL U2205 ( .A0(n3148), .A1(n3188), .B0(n3189), .B1(n290), .Y(n1971) );
  OAI22XL U2206 ( .A0(n3146), .A1(n3188), .B0(n3189), .B1(n289), .Y(n1972) );
  OAI22XL U2207 ( .A0(n3144), .A1(n3191), .B0(n3189), .B1(n288), .Y(n1973) );
  OAI22XL U2208 ( .A0(n3142), .A1(n3191), .B0(n3189), .B1(n287), .Y(n1974) );
  OAI22XL U2209 ( .A0(n3140), .A1(n112), .B0(n3190), .B1(n286), .Y(n1975) );
  OAI22XL U2210 ( .A0(n3138), .A1(n112), .B0(n3190), .B1(n285), .Y(n1976) );
  OAI22XL U2211 ( .A0(n3136), .A1(n3188), .B0(n3190), .B1(n284), .Y(n1977) );
  OAI22XL U2212 ( .A0(n3134), .A1(n3188), .B0(n3190), .B1(n283), .Y(n1978) );
  OAI22XL U2213 ( .A0(n3132), .A1(n3188), .B0(n3190), .B1(n282), .Y(n1979) );
  OAI22XL U2214 ( .A0(n3130), .A1(n3188), .B0(n3190), .B1(n281), .Y(n1980) );
  OAI22XL U2215 ( .A0(n3128), .A1(n112), .B0(n3190), .B1(n280), .Y(n1981) );
  OAI22XL U2216 ( .A0(n3126), .A1(n112), .B0(n3190), .B1(n279), .Y(n1982) );
  OAI22XL U2217 ( .A0(n3124), .A1(n3188), .B0(n3190), .B1(n278), .Y(n1983) );
  OAI22XL U2218 ( .A0(n3122), .A1(n3188), .B0(n3190), .B1(n277), .Y(n1984) );
  OAI22XL U2219 ( .A0(n3120), .A1(n3188), .B0(n3190), .B1(n276), .Y(n1985) );
  OAI22XL U2220 ( .A0(n3118), .A1(n3188), .B0(n3190), .B1(n275), .Y(n1986) );
  OAI22XL U2221 ( .A0(n3164), .A1(n3187), .B0(n3185), .B1(n266), .Y(n1995) );
  OAI22XL U2222 ( .A0(n3162), .A1(n3187), .B0(n3185), .B1(n265), .Y(n1996) );
  OAI22XL U2223 ( .A0(n3160), .A1(n3187), .B0(n3185), .B1(n264), .Y(n1997) );
  OAI22XL U2224 ( .A0(n3158), .A1(n3187), .B0(n3185), .B1(n263), .Y(n1998) );
  OAI22XL U2225 ( .A0(n3156), .A1(n3184), .B0(n3185), .B1(n262), .Y(n1999) );
  OAI22XL U2226 ( .A0(n3154), .A1(n3187), .B0(n3185), .B1(n261), .Y(n2000) );
  OAI22XL U2227 ( .A0(n3152), .A1(n3184), .B0(n3185), .B1(n260), .Y(n2001) );
  OAI22XL U2228 ( .A0(n3150), .A1(n3184), .B0(n3185), .B1(n259), .Y(n2002) );
  OAI22XL U2229 ( .A0(n3148), .A1(n3187), .B0(n3185), .B1(n258), .Y(n2003) );
  OAI22XL U2230 ( .A0(n3146), .A1(n3187), .B0(n3185), .B1(n257), .Y(n2004) );
  OAI22XL U2231 ( .A0(n3144), .A1(n3184), .B0(n3185), .B1(n256), .Y(n2005) );
  OAI22XL U2232 ( .A0(n3142), .A1(n3187), .B0(n3185), .B1(n255), .Y(n2006) );
  OAI22XL U2233 ( .A0(n3140), .A1(n3184), .B0(n3186), .B1(n254), .Y(n2007) );
  OAI22XL U2234 ( .A0(n3138), .A1(n3184), .B0(n3186), .B1(n253), .Y(n2008) );
  OAI22XL U2235 ( .A0(n3136), .A1(n3184), .B0(n3186), .B1(n252), .Y(n2009) );
  OAI22XL U2236 ( .A0(n3134), .A1(n3184), .B0(n3186), .B1(n251), .Y(n2010) );
  OAI22XL U2237 ( .A0(n3132), .A1(n115), .B0(n3186), .B1(n250), .Y(n2011) );
  OAI22XL U2238 ( .A0(n3130), .A1(n115), .B0(n3186), .B1(n249), .Y(n2012) );
  OAI22XL U2239 ( .A0(n3128), .A1(n115), .B0(n3186), .B1(n248), .Y(n2013) );
  OAI22XL U2240 ( .A0(n3126), .A1(n115), .B0(n3186), .B1(n247), .Y(n2014) );
  OAI22XL U2241 ( .A0(n3124), .A1(n115), .B0(n3186), .B1(n246), .Y(n2015) );
  OAI22XL U2242 ( .A0(n3122), .A1(n3184), .B0(n3186), .B1(n245), .Y(n2016) );
  OAI22XL U2243 ( .A0(n3120), .A1(n3184), .B0(n3186), .B1(n244), .Y(n2017) );
  OAI22XL U2244 ( .A0(n3118), .A1(n3184), .B0(n3186), .B1(n243), .Y(n2018) );
  OAI22XL U2245 ( .A0(n3164), .A1(n3183), .B0(n3181), .B1(n234), .Y(n2027) );
  OAI22XL U2246 ( .A0(n3162), .A1(n3183), .B0(n3181), .B1(n233), .Y(n2028) );
  OAI22XL U2247 ( .A0(n3160), .A1(n3183), .B0(n3181), .B1(n232), .Y(n2029) );
  OAI22XL U2248 ( .A0(n3158), .A1(n3183), .B0(n3181), .B1(n231), .Y(n2030) );
  OAI22XL U2249 ( .A0(n3156), .A1(n3180), .B0(n3181), .B1(n230), .Y(n2031) );
  OAI22XL U2250 ( .A0(n3154), .A1(n3180), .B0(n3181), .B1(n229), .Y(n2032) );
  OAI22XL U2251 ( .A0(n3152), .A1(n3180), .B0(n3181), .B1(n228), .Y(n2033) );
  OAI22XL U2252 ( .A0(n3150), .A1(n3180), .B0(n3181), .B1(n227), .Y(n2034) );
  OAI22XL U2253 ( .A0(n3148), .A1(n3180), .B0(n3181), .B1(n226), .Y(n2035) );
  OAI22XL U2254 ( .A0(n3146), .A1(n3180), .B0(n3181), .B1(n225), .Y(n2036) );
  OAI22XL U2255 ( .A0(n3144), .A1(n3183), .B0(n3181), .B1(n224), .Y(n2037) );
  OAI22XL U2256 ( .A0(n3142), .A1(n3183), .B0(n3181), .B1(n223), .Y(n2038) );
  OAI22XL U2257 ( .A0(n3140), .A1(n117), .B0(n3182), .B1(n222), .Y(n2039) );
  OAI22XL U2258 ( .A0(n3138), .A1(n117), .B0(n3182), .B1(n221), .Y(n2040) );
  OAI22XL U2259 ( .A0(n3136), .A1(n3180), .B0(n3182), .B1(n220), .Y(n2041) );
  OAI22XL U2260 ( .A0(n3134), .A1(n3180), .B0(n3182), .B1(n219), .Y(n2042) );
  OAI22XL U2261 ( .A0(n3132), .A1(n3180), .B0(n3182), .B1(n218), .Y(n2043) );
  OAI22XL U2262 ( .A0(n3130), .A1(n3180), .B0(n3182), .B1(n217), .Y(n2044) );
  OAI22XL U2263 ( .A0(n3128), .A1(n117), .B0(n3182), .B1(n216), .Y(n2045) );
  OAI22XL U2264 ( .A0(n3126), .A1(n117), .B0(n3182), .B1(n215), .Y(n2046) );
  OAI22XL U2265 ( .A0(n3124), .A1(n3180), .B0(n3182), .B1(n214), .Y(n2047) );
  OAI22XL U2266 ( .A0(n3122), .A1(n3180), .B0(n3182), .B1(n213), .Y(n2048) );
  OAI22XL U2267 ( .A0(n3120), .A1(n3180), .B0(n3182), .B1(n212), .Y(n2049) );
  OAI22XL U2268 ( .A0(n3118), .A1(n3180), .B0(n3182), .B1(n211), .Y(n2050) );
  OAI22XL U2269 ( .A0(n3164), .A1(n3179), .B0(n3177), .B1(n202), .Y(n2059) );
  OAI22XL U2270 ( .A0(n3162), .A1(n3179), .B0(n3177), .B1(n201), .Y(n2060) );
  OAI22XL U2271 ( .A0(n3160), .A1(n3179), .B0(n3177), .B1(n200), .Y(n2061) );
  OAI22XL U2272 ( .A0(n3158), .A1(n3179), .B0(n3177), .B1(n199), .Y(n2062) );
  OAI22XL U2273 ( .A0(n3156), .A1(n3176), .B0(n3177), .B1(n198), .Y(n2063) );
  OAI22XL U2274 ( .A0(n3154), .A1(n3179), .B0(n3177), .B1(n197), .Y(n2064) );
  OAI22XL U2275 ( .A0(n3152), .A1(n3176), .B0(n3177), .B1(n196), .Y(n2065) );
  OAI22XL U2276 ( .A0(n3150), .A1(n3176), .B0(n3177), .B1(n195), .Y(n2066) );
  OAI22XL U2277 ( .A0(n3148), .A1(n3179), .B0(n3177), .B1(n194), .Y(n2067) );
  OAI22XL U2278 ( .A0(n3146), .A1(n3179), .B0(n3177), .B1(n193), .Y(n2068) );
  OAI22XL U2279 ( .A0(n3144), .A1(n3176), .B0(n3177), .B1(n192), .Y(n2069) );
  OAI22XL U2280 ( .A0(n3142), .A1(n3179), .B0(n3177), .B1(n191), .Y(n2070) );
  OAI22XL U2281 ( .A0(n3140), .A1(n3176), .B0(n3178), .B1(n190), .Y(n2071) );
  OAI22XL U2282 ( .A0(n3138), .A1(n3176), .B0(n3178), .B1(n189), .Y(n2072) );
  OAI22XL U2283 ( .A0(n3136), .A1(n3176), .B0(n3178), .B1(n188), .Y(n2073) );
  OAI22XL U2284 ( .A0(n3134), .A1(n3176), .B0(n3178), .B1(n187), .Y(n2074) );
  OAI22XL U2285 ( .A0(n3132), .A1(n120), .B0(n3178), .B1(n186), .Y(n2075) );
  OAI22XL U2286 ( .A0(n3130), .A1(n120), .B0(n3178), .B1(n185), .Y(n2076) );
  OAI22XL U2287 ( .A0(n3128), .A1(n120), .B0(n3178), .B1(n184), .Y(n2077) );
  OAI22XL U2288 ( .A0(n3126), .A1(n120), .B0(n3178), .B1(n183), .Y(n2078) );
  OAI22XL U2289 ( .A0(n3124), .A1(n120), .B0(n3178), .B1(n182), .Y(n2079) );
  OAI22XL U2290 ( .A0(n3122), .A1(n3176), .B0(n3178), .B1(n181), .Y(n2080) );
  OAI22XL U2291 ( .A0(n3120), .A1(n3176), .B0(n3178), .B1(n180), .Y(n2081) );
  OAI22XL U2292 ( .A0(n3118), .A1(n3176), .B0(n3178), .B1(n179), .Y(n2082) );
  OAI22XL U2293 ( .A0(n3164), .A1(n3175), .B0(n3173), .B1(n170), .Y(n2091) );
  OAI22XL U2294 ( .A0(n3162), .A1(n3175), .B0(n3173), .B1(n169), .Y(n2092) );
  OAI22XL U2295 ( .A0(n3160), .A1(n3175), .B0(n3173), .B1(n168), .Y(n2093) );
  OAI22XL U2296 ( .A0(n3158), .A1(n3175), .B0(n3173), .B1(n167), .Y(n2094) );
  OAI22XL U2297 ( .A0(n3156), .A1(n3172), .B0(n3173), .B1(n166), .Y(n2095) );
  OAI22XL U2298 ( .A0(n3154), .A1(n3172), .B0(n3173), .B1(n165), .Y(n2096) );
  OAI22XL U2299 ( .A0(n3152), .A1(n3172), .B0(n3173), .B1(n164), .Y(n2097) );
  OAI22XL U2300 ( .A0(n3150), .A1(n3172), .B0(n3173), .B1(n163), .Y(n2098) );
  OAI22XL U2301 ( .A0(n3148), .A1(n3172), .B0(n3173), .B1(n162), .Y(n2099) );
  OAI22XL U2302 ( .A0(n3146), .A1(n3172), .B0(n3173), .B1(n161), .Y(n2100) );
  OAI22XL U2303 ( .A0(n3144), .A1(n3175), .B0(n3173), .B1(n160), .Y(n2101) );
  OAI22XL U2304 ( .A0(n3142), .A1(n3175), .B0(n3173), .B1(n159), .Y(n2102) );
  OAI22XL U2305 ( .A0(n3140), .A1(n123), .B0(n3174), .B1(n158), .Y(n2103) );
  OAI22XL U2306 ( .A0(n3138), .A1(n123), .B0(n3174), .B1(n157), .Y(n2104) );
  OAI22XL U2307 ( .A0(n3136), .A1(n3172), .B0(n3174), .B1(n156), .Y(n2105) );
  OAI22XL U2308 ( .A0(n3134), .A1(n3172), .B0(n3174), .B1(n155), .Y(n2106) );
  OAI22XL U2309 ( .A0(n3132), .A1(n3172), .B0(n3174), .B1(n154), .Y(n2107) );
  OAI22XL U2310 ( .A0(n3130), .A1(n3172), .B0(n3174), .B1(n153), .Y(n2108) );
  OAI22XL U2311 ( .A0(n3128), .A1(n123), .B0(n3174), .B1(n152), .Y(n2109) );
  OAI22XL U2312 ( .A0(n3126), .A1(n123), .B0(n3174), .B1(n151), .Y(n2110) );
  OAI22XL U2313 ( .A0(n3124), .A1(n3172), .B0(n3174), .B1(n150), .Y(n2111) );
  OAI22XL U2314 ( .A0(n3122), .A1(n3172), .B0(n3174), .B1(n149), .Y(n2112) );
  OAI22XL U2315 ( .A0(n3120), .A1(n3172), .B0(n3174), .B1(n148), .Y(n2113) );
  OAI22XL U2316 ( .A0(n3118), .A1(n3172), .B0(n3174), .B1(n147), .Y(n2114) );
  OAI22XL U2317 ( .A0(n3292), .A1(n3165), .B0(n3294), .B1(n1130), .Y(n1131) );
  OAI22XL U2318 ( .A0(n3293), .A1(n3163), .B0(n3294), .B1(n1129), .Y(n1132) );
  OAI22XL U2319 ( .A0(n3292), .A1(n3161), .B0(n3294), .B1(n1128), .Y(n1133) );
  OAI22XL U2320 ( .A0(n3292), .A1(n3159), .B0(n3294), .B1(n1127), .Y(n1134) );
  OAI22XL U2321 ( .A0(n3292), .A1(n3157), .B0(n3294), .B1(n1126), .Y(n1135) );
  OAI22XL U2322 ( .A0(n3292), .A1(n3155), .B0(n3294), .B1(n1125), .Y(n1136) );
  OAI22XL U2323 ( .A0(n9), .A1(n3153), .B0(n3294), .B1(n1124), .Y(n1137) );
  OAI22XL U2324 ( .A0(n9), .A1(n3151), .B0(n3295), .B1(n1123), .Y(n1138) );
  OAI22XL U2325 ( .A0(n9), .A1(n3149), .B0(n3295), .B1(n1122), .Y(n1139) );
  OAI22XL U2326 ( .A0(n9), .A1(n3147), .B0(n3295), .B1(n1121), .Y(n1140) );
  OAI22XL U2327 ( .A0(n9), .A1(n3145), .B0(n3295), .B1(n1120), .Y(n1141) );
  OAI22XL U2328 ( .A0(n9), .A1(n3143), .B0(n3295), .B1(n1119), .Y(n1142) );
  OAI22XL U2329 ( .A0(n3292), .A1(n3141), .B0(n3294), .B1(n1118), .Y(n1143) );
  OAI22XL U2330 ( .A0(n3292), .A1(n3139), .B0(n3294), .B1(n1117), .Y(n1144) );
  OAI22XL U2331 ( .A0(n3292), .A1(n3137), .B0(n3295), .B1(n1116), .Y(n1145) );
  OAI22XL U2332 ( .A0(n3292), .A1(n3135), .B0(n3294), .B1(n1115), .Y(n1146) );
  OAI22XL U2333 ( .A0(n3292), .A1(n3133), .B0(n3295), .B1(n1114), .Y(n1147) );
  OAI22XL U2334 ( .A0(n3292), .A1(n3131), .B0(n3294), .B1(n1113), .Y(n1148) );
  OAI22XL U2335 ( .A0(n3292), .A1(n3129), .B0(n3295), .B1(n1112), .Y(n1149) );
  OAI22XL U2336 ( .A0(n3292), .A1(n3127), .B0(n3294), .B1(n1111), .Y(n1150) );
  OAI22XL U2337 ( .A0(n3292), .A1(n3125), .B0(n3295), .B1(n1110), .Y(n1151) );
  OAI22XL U2338 ( .A0(n3292), .A1(n3123), .B0(n3295), .B1(n1109), .Y(n1152) );
  OAI22XL U2339 ( .A0(n3292), .A1(n3121), .B0(n3295), .B1(n1108), .Y(n1153) );
  OAI22XL U2340 ( .A0(n3292), .A1(n3119), .B0(n3295), .B1(n1107), .Y(n1154) );
  OAI22XL U2341 ( .A0(n3293), .A1(n3117), .B0(n3295), .B1(n1106), .Y(n1155) );
  OAI22XL U2342 ( .A0(n3293), .A1(n3115), .B0(n3294), .B1(n1105), .Y(n1156) );
  OAI22XL U2343 ( .A0(n3293), .A1(n3113), .B0(n3294), .B1(n1104), .Y(n1157) );
  OAI22XL U2344 ( .A0(n3293), .A1(n3111), .B0(n3295), .B1(n1103), .Y(n1158) );
  OAI22XL U2345 ( .A0(n3293), .A1(n3109), .B0(n3294), .B1(n1102), .Y(n1159) );
  OAI22XL U2346 ( .A0(n3293), .A1(n3107), .B0(n3295), .B1(n1101), .Y(n1160) );
  OAI22XL U2347 ( .A0(n3293), .A1(n3105), .B0(n3294), .B1(n1100), .Y(n1161) );
  OAI22XL U2348 ( .A0(n3293), .A1(n3103), .B0(n3295), .B1(n1099), .Y(n1162) );
  OAI22XL U2349 ( .A0(n3117), .A1(n3284), .B0(n3286), .B1(n1042), .Y(n1219) );
  OAI22XL U2350 ( .A0(n3115), .A1(n49), .B0(n3286), .B1(n1041), .Y(n1220) );
  OAI22XL U2351 ( .A0(n3113), .A1(n49), .B0(n3286), .B1(n1040), .Y(n1221) );
  OAI22XL U2352 ( .A0(n3111), .A1(n3284), .B0(n3286), .B1(n1039), .Y(n1222) );
  OAI22XL U2353 ( .A0(n3109), .A1(n3284), .B0(n3286), .B1(n1038), .Y(n1223) );
  OAI22XL U2354 ( .A0(n3107), .A1(n3284), .B0(n3286), .B1(n1037), .Y(n1224) );
  OAI22XL U2355 ( .A0(n3105), .A1(n3287), .B0(n3286), .B1(n1036), .Y(n1225) );
  OAI22XL U2356 ( .A0(n3103), .A1(n3284), .B0(n3286), .B1(n1035), .Y(n1226) );
  OAI22XL U2357 ( .A0(n3117), .A1(n3283), .B0(n3281), .B1(n1010), .Y(n1251) );
  OAI22XL U2358 ( .A0(n3115), .A1(n3283), .B0(n3282), .B1(n1009), .Y(n1252) );
  OAI22XL U2359 ( .A0(n3113), .A1(n3283), .B0(n3281), .B1(n1008), .Y(n1253) );
  OAI22XL U2360 ( .A0(n3111), .A1(n3283), .B0(n3282), .B1(n1007), .Y(n1254) );
  OAI22XL U2361 ( .A0(n3109), .A1(n3280), .B0(n3281), .B1(n1006), .Y(n1255) );
  OAI22XL U2362 ( .A0(n3107), .A1(n3280), .B0(n3282), .B1(n1005), .Y(n1256) );
  OAI22XL U2363 ( .A0(n3105), .A1(n3283), .B0(n3281), .B1(n1004), .Y(n1257) );
  OAI22XL U2364 ( .A0(n3103), .A1(n3280), .B0(n3282), .B1(n1003), .Y(n1258) );
  OAI22XL U2365 ( .A0(n3117), .A1(n3276), .B0(n3277), .B1(n978), .Y(n1283) );
  OAI22XL U2366 ( .A0(n3115), .A1(n54), .B0(n3278), .B1(n977), .Y(n1284) );
  OAI22XL U2367 ( .A0(n3113), .A1(n54), .B0(n3277), .B1(n976), .Y(n1285) );
  OAI22XL U2368 ( .A0(n3111), .A1(n3276), .B0(n3278), .B1(n975), .Y(n1286) );
  OAI22XL U2369 ( .A0(n3109), .A1(n3276), .B0(n3277), .B1(n974), .Y(n1287) );
  OAI22XL U2370 ( .A0(n3107), .A1(n3276), .B0(n3278), .B1(n973), .Y(n1288) );
  OAI22XL U2371 ( .A0(n3105), .A1(n3279), .B0(n3277), .B1(n972), .Y(n1289) );
  OAI22XL U2372 ( .A0(n3103), .A1(n3276), .B0(n3278), .B1(n971), .Y(n1290) );
  OAI22XL U2373 ( .A0(n3117), .A1(n3275), .B0(n3273), .B1(n946), .Y(n1315) );
  OAI22XL U2374 ( .A0(n3115), .A1(n3275), .B0(n3274), .B1(n945), .Y(n1316) );
  OAI22XL U2375 ( .A0(n3113), .A1(n3275), .B0(n3273), .B1(n944), .Y(n1317) );
  OAI22XL U2376 ( .A0(n3111), .A1(n3275), .B0(n3274), .B1(n943), .Y(n1318) );
  OAI22XL U2377 ( .A0(n3109), .A1(n3272), .B0(n3273), .B1(n942), .Y(n1319) );
  OAI22XL U2378 ( .A0(n3107), .A1(n3272), .B0(n3274), .B1(n941), .Y(n1320) );
  OAI22XL U2379 ( .A0(n3105), .A1(n3275), .B0(n3273), .B1(n940), .Y(n1321) );
  OAI22XL U2380 ( .A0(n3103), .A1(n3272), .B0(n3274), .B1(n939), .Y(n1322) );
  OAI22XL U2381 ( .A0(n3117), .A1(n3268), .B0(n3269), .B1(n914), .Y(n1347) );
  OAI22XL U2382 ( .A0(n3115), .A1(n60), .B0(n3270), .B1(n913), .Y(n1348) );
  OAI22XL U2383 ( .A0(n3113), .A1(n60), .B0(n3269), .B1(n912), .Y(n1349) );
  OAI22XL U2384 ( .A0(n3111), .A1(n3268), .B0(n3270), .B1(n911), .Y(n1350) );
  OAI22XL U2385 ( .A0(n3109), .A1(n3268), .B0(n3269), .B1(n910), .Y(n1351) );
  OAI22XL U2386 ( .A0(n3107), .A1(n3268), .B0(n3270), .B1(n909), .Y(n1352) );
  OAI22XL U2387 ( .A0(n3105), .A1(n3271), .B0(n3269), .B1(n908), .Y(n1353) );
  OAI22XL U2388 ( .A0(n3103), .A1(n3268), .B0(n3270), .B1(n907), .Y(n1354) );
  OAI22XL U2389 ( .A0(n3117), .A1(n3264), .B0(n3265), .B1(n882), .Y(n1379) );
  OAI22XL U2390 ( .A0(n3115), .A1(n3264), .B0(n3266), .B1(n881), .Y(n1380) );
  OAI22XL U2391 ( .A0(n3113), .A1(n3264), .B0(n3265), .B1(n880), .Y(n1381) );
  OAI22XL U2392 ( .A0(n3111), .A1(n64), .B0(n3266), .B1(n879), .Y(n1382) );
  OAI22XL U2393 ( .A0(n3109), .A1(n3264), .B0(n3265), .B1(n878), .Y(n1383) );
  OAI22XL U2394 ( .A0(n3107), .A1(n3267), .B0(n3266), .B1(n877), .Y(n1384) );
  OAI22XL U2395 ( .A0(n3105), .A1(n3267), .B0(n3265), .B1(n876), .Y(n1385) );
  OAI22XL U2396 ( .A0(n3103), .A1(n3264), .B0(n3266), .B1(n875), .Y(n1386) );
  OAI22XL U2397 ( .A0(n3117), .A1(n3260), .B0(n3261), .B1(n850), .Y(n1411) );
  OAI22XL U2398 ( .A0(n3115), .A1(n3260), .B0(n3262), .B1(n849), .Y(n1412) );
  OAI22XL U2399 ( .A0(n3113), .A1(n3260), .B0(n3261), .B1(n848), .Y(n1413) );
  OAI22XL U2400 ( .A0(n3111), .A1(n67), .B0(n3262), .B1(n847), .Y(n1414) );
  OAI22XL U2401 ( .A0(n3109), .A1(n3260), .B0(n3261), .B1(n846), .Y(n1415) );
  OAI22XL U2402 ( .A0(n3107), .A1(n3263), .B0(n3262), .B1(n845), .Y(n1416) );
  OAI22XL U2403 ( .A0(n3105), .A1(n3263), .B0(n3261), .B1(n844), .Y(n1417) );
  OAI22XL U2404 ( .A0(n3103), .A1(n3260), .B0(n3262), .B1(n843), .Y(n1418) );
  OAI22XL U2405 ( .A0(n3117), .A1(n3256), .B0(n3257), .B1(n818), .Y(n1443) );
  OAI22XL U2406 ( .A0(n3115), .A1(n3256), .B0(n3258), .B1(n817), .Y(n1444) );
  OAI22XL U2407 ( .A0(n3113), .A1(n3256), .B0(n3257), .B1(n816), .Y(n1445) );
  OAI22XL U2408 ( .A0(n3111), .A1(n70), .B0(n3258), .B1(n815), .Y(n1446) );
  OAI22XL U2409 ( .A0(n3109), .A1(n3256), .B0(n3257), .B1(n814), .Y(n1447) );
  OAI22XL U2410 ( .A0(n3107), .A1(n3259), .B0(n3258), .B1(n813), .Y(n1448) );
  OAI22XL U2411 ( .A0(n3105), .A1(n3259), .B0(n3257), .B1(n812), .Y(n1449) );
  OAI22XL U2412 ( .A0(n3103), .A1(n3256), .B0(n3258), .B1(n811), .Y(n1450) );
  OAI22XL U2413 ( .A0(n3117), .A1(n3252), .B0(n3253), .B1(n786), .Y(n1475) );
  OAI22XL U2414 ( .A0(n3115), .A1(n3252), .B0(n3254), .B1(n785), .Y(n1476) );
  OAI22XL U2415 ( .A0(n3113), .A1(n3252), .B0(n3253), .B1(n784), .Y(n1477) );
  OAI22XL U2416 ( .A0(n3111), .A1(n72), .B0(n3254), .B1(n783), .Y(n1478) );
  OAI22XL U2417 ( .A0(n3109), .A1(n3252), .B0(n3253), .B1(n782), .Y(n1479) );
  OAI22XL U2418 ( .A0(n3107), .A1(n3255), .B0(n3254), .B1(n781), .Y(n1480) );
  OAI22XL U2419 ( .A0(n3105), .A1(n3255), .B0(n3253), .B1(n780), .Y(n1481) );
  OAI22XL U2420 ( .A0(n3103), .A1(n3252), .B0(n3254), .B1(n779), .Y(n1482) );
  OAI22XL U2421 ( .A0(n3117), .A1(n3248), .B0(n3249), .B1(n754), .Y(n1507) );
  OAI22XL U2422 ( .A0(n3115), .A1(n3248), .B0(n3250), .B1(n753), .Y(n1508) );
  OAI22XL U2423 ( .A0(n3113), .A1(n3248), .B0(n3249), .B1(n752), .Y(n1509) );
  OAI22XL U2424 ( .A0(n3111), .A1(n74), .B0(n3250), .B1(n751), .Y(n1510) );
  OAI22XL U2425 ( .A0(n3109), .A1(n3248), .B0(n3249), .B1(n750), .Y(n1511) );
  OAI22XL U2426 ( .A0(n3107), .A1(n3251), .B0(n3250), .B1(n749), .Y(n1512) );
  OAI22XL U2427 ( .A0(n3105), .A1(n3251), .B0(n3249), .B1(n748), .Y(n1513) );
  OAI22XL U2428 ( .A0(n3103), .A1(n3248), .B0(n3250), .B1(n747), .Y(n1514) );
  OAI22XL U2429 ( .A0(n3117), .A1(n3244), .B0(n3245), .B1(n722), .Y(n1539) );
  OAI22XL U2430 ( .A0(n3115), .A1(n3244), .B0(n3246), .B1(n721), .Y(n1540) );
  OAI22XL U2431 ( .A0(n3113), .A1(n3244), .B0(n3245), .B1(n720), .Y(n1541) );
  OAI22XL U2432 ( .A0(n3111), .A1(n76), .B0(n3246), .B1(n719), .Y(n1542) );
  OAI22XL U2433 ( .A0(n3109), .A1(n3244), .B0(n3245), .B1(n718), .Y(n1543) );
  OAI22XL U2434 ( .A0(n3107), .A1(n3247), .B0(n3246), .B1(n717), .Y(n1544) );
  OAI22XL U2435 ( .A0(n3105), .A1(n3247), .B0(n3245), .B1(n716), .Y(n1545) );
  OAI22XL U2436 ( .A0(n3103), .A1(n3244), .B0(n3246), .B1(n715), .Y(n1546) );
  OAI22XL U2437 ( .A0(n3117), .A1(n3240), .B0(n3241), .B1(n690), .Y(n1571) );
  OAI22XL U2438 ( .A0(n3115), .A1(n3240), .B0(n3242), .B1(n689), .Y(n1572) );
  OAI22XL U2439 ( .A0(n3113), .A1(n3240), .B0(n3241), .B1(n688), .Y(n1573) );
  OAI22XL U2440 ( .A0(n3111), .A1(n78), .B0(n3242), .B1(n687), .Y(n1574) );
  OAI22XL U2441 ( .A0(n3109), .A1(n3240), .B0(n3241), .B1(n686), .Y(n1575) );
  OAI22XL U2442 ( .A0(n3107), .A1(n3243), .B0(n3242), .B1(n685), .Y(n1576) );
  OAI22XL U2443 ( .A0(n3105), .A1(n3243), .B0(n3241), .B1(n684), .Y(n1577) );
  OAI22XL U2444 ( .A0(n3103), .A1(n3240), .B0(n3242), .B1(n683), .Y(n1578) );
  OAI22XL U2445 ( .A0(n3117), .A1(n3236), .B0(n3237), .B1(n658), .Y(n1603) );
  OAI22XL U2446 ( .A0(n3115), .A1(n3236), .B0(n3238), .B1(n657), .Y(n1604) );
  OAI22XL U2447 ( .A0(n3113), .A1(n3236), .B0(n3237), .B1(n656), .Y(n1605) );
  OAI22XL U2448 ( .A0(n3111), .A1(n81), .B0(n3238), .B1(n655), .Y(n1606) );
  OAI22XL U2449 ( .A0(n3109), .A1(n3236), .B0(n3237), .B1(n654), .Y(n1607) );
  OAI22XL U2450 ( .A0(n3107), .A1(n3239), .B0(n3238), .B1(n653), .Y(n1608) );
  OAI22XL U2451 ( .A0(n3105), .A1(n3239), .B0(n3237), .B1(n652), .Y(n1609) );
  OAI22XL U2452 ( .A0(n3103), .A1(n3236), .B0(n3238), .B1(n651), .Y(n1610) );
  OAI22XL U2453 ( .A0(n3117), .A1(n3235), .B0(n3233), .B1(n626), .Y(n1635) );
  OAI22XL U2454 ( .A0(n3115), .A1(n3235), .B0(n3233), .B1(n625), .Y(n1636) );
  OAI22XL U2455 ( .A0(n3113), .A1(n3235), .B0(n3233), .B1(n624), .Y(n1637) );
  OAI22XL U2456 ( .A0(n3111), .A1(n3235), .B0(n3233), .B1(n623), .Y(n1638) );
  OAI22XL U2457 ( .A0(n3109), .A1(n3232), .B0(n3233), .B1(n622), .Y(n1639) );
  OAI22XL U2458 ( .A0(n3107), .A1(n3232), .B0(n3233), .B1(n621), .Y(n1640) );
  OAI22XL U2459 ( .A0(n3105), .A1(n3232), .B0(n3233), .B1(n620), .Y(n1641) );
  OAI22XL U2460 ( .A0(n3103), .A1(n3235), .B0(n3233), .B1(n619), .Y(n1642) );
  OAI22XL U2461 ( .A0(n3117), .A1(n3231), .B0(n3229), .B1(n594), .Y(n1667) );
  OAI22XL U2462 ( .A0(n3115), .A1(n3231), .B0(n3229), .B1(n593), .Y(n1668) );
  OAI22XL U2463 ( .A0(n3113), .A1(n3231), .B0(n3229), .B1(n592), .Y(n1669) );
  OAI22XL U2464 ( .A0(n3111), .A1(n3231), .B0(n3229), .B1(n591), .Y(n1670) );
  OAI22XL U2465 ( .A0(n3109), .A1(n3228), .B0(n3229), .B1(n590), .Y(n1671) );
  OAI22XL U2466 ( .A0(n3107), .A1(n3228), .B0(n3229), .B1(n589), .Y(n1672) );
  OAI22XL U2467 ( .A0(n3105), .A1(n3228), .B0(n3229), .B1(n588), .Y(n1673) );
  OAI22XL U2468 ( .A0(n3103), .A1(n3231), .B0(n3229), .B1(n587), .Y(n1674) );
  OAI22XL U2469 ( .A0(n3117), .A1(n3227), .B0(n3225), .B1(n562), .Y(n1699) );
  OAI22XL U2470 ( .A0(n3115), .A1(n3227), .B0(n3225), .B1(n561), .Y(n1700) );
  OAI22XL U2471 ( .A0(n3113), .A1(n3227), .B0(n3225), .B1(n560), .Y(n1701) );
  OAI22XL U2472 ( .A0(n3111), .A1(n3227), .B0(n3225), .B1(n559), .Y(n1702) );
  OAI22XL U2473 ( .A0(n3109), .A1(n3224), .B0(n3225), .B1(n558), .Y(n1703) );
  OAI22XL U2474 ( .A0(n3107), .A1(n3224), .B0(n3225), .B1(n557), .Y(n1704) );
  OAI22XL U2475 ( .A0(n3105), .A1(n3224), .B0(n3225), .B1(n556), .Y(n1705) );
  OAI22XL U2476 ( .A0(n3103), .A1(n3227), .B0(n3225), .B1(n555), .Y(n1706) );
  OAI22XL U2477 ( .A0(n3117), .A1(n3223), .B0(n3221), .B1(n530), .Y(n1731) );
  OAI22XL U2478 ( .A0(n3115), .A1(n3223), .B0(n3221), .B1(n529), .Y(n1732) );
  OAI22XL U2479 ( .A0(n3113), .A1(n3223), .B0(n3221), .B1(n528), .Y(n1733) );
  OAI22XL U2480 ( .A0(n3111), .A1(n3223), .B0(n3221), .B1(n527), .Y(n1734) );
  OAI22XL U2481 ( .A0(n3109), .A1(n3220), .B0(n3221), .B1(n526), .Y(n1735) );
  OAI22XL U2482 ( .A0(n3107), .A1(n3220), .B0(n3221), .B1(n525), .Y(n1736) );
  OAI22XL U2483 ( .A0(n3105), .A1(n3220), .B0(n3221), .B1(n524), .Y(n1737) );
  OAI22XL U2484 ( .A0(n3103), .A1(n3223), .B0(n3221), .B1(n523), .Y(n1738) );
  OAI22XL U2485 ( .A0(n3117), .A1(n94), .B0(n3218), .B1(n498), .Y(n1763) );
  OAI22XL U2486 ( .A0(n3115), .A1(n94), .B0(n3218), .B1(n497), .Y(n1764) );
  OAI22XL U2487 ( .A0(n3113), .A1(n3216), .B0(n3218), .B1(n496), .Y(n1765) );
  OAI22XL U2488 ( .A0(n3111), .A1(n3216), .B0(n3218), .B1(n495), .Y(n1766) );
  OAI22XL U2489 ( .A0(n3109), .A1(n94), .B0(n3218), .B1(n494), .Y(n1767) );
  OAI22XL U2490 ( .A0(n3107), .A1(n3219), .B0(n3218), .B1(n493), .Y(n1768) );
  OAI22XL U2491 ( .A0(n3105), .A1(n3216), .B0(n3218), .B1(n492), .Y(n1769) );
  OAI22XL U2492 ( .A0(n3103), .A1(n94), .B0(n3218), .B1(n491), .Y(n1770) );
  OAI22XL U2493 ( .A0(n3116), .A1(n3212), .B0(n3214), .B1(n466), .Y(n1795) );
  OAI22XL U2494 ( .A0(n3114), .A1(n3212), .B0(n3215), .B1(n465), .Y(n1796) );
  OAI22XL U2495 ( .A0(n3112), .A1(n3212), .B0(n3214), .B1(n464), .Y(n1797) );
  OAI22XL U2496 ( .A0(n3110), .A1(n3213), .B0(n3215), .B1(n463), .Y(n1798) );
  OAI22XL U2497 ( .A0(n3108), .A1(n3213), .B0(n3214), .B1(n462), .Y(n1799) );
  OAI22XL U2498 ( .A0(n3106), .A1(n3212), .B0(n3215), .B1(n461), .Y(n1800) );
  OAI22XL U2499 ( .A0(n3104), .A1(n3213), .B0(n3214), .B1(n460), .Y(n1801) );
  OAI22XL U2500 ( .A0(n3102), .A1(n3213), .B0(n3215), .B1(n459), .Y(n1802) );
  OAI22XL U2501 ( .A0(n3116), .A1(n3208), .B0(n3210), .B1(n434), .Y(n1827) );
  OAI22XL U2502 ( .A0(n3114), .A1(n3208), .B0(n3211), .B1(n433), .Y(n1828) );
  OAI22XL U2503 ( .A0(n3112), .A1(n3208), .B0(n3210), .B1(n432), .Y(n1829) );
  OAI22XL U2504 ( .A0(n3110), .A1(n3209), .B0(n3211), .B1(n431), .Y(n1830) );
  OAI22XL U2505 ( .A0(n3108), .A1(n3209), .B0(n3210), .B1(n430), .Y(n1831) );
  OAI22XL U2506 ( .A0(n3106), .A1(n3208), .B0(n3211), .B1(n429), .Y(n1832) );
  OAI22XL U2507 ( .A0(n3104), .A1(n3209), .B0(n3210), .B1(n428), .Y(n1833) );
  OAI22XL U2508 ( .A0(n3102), .A1(n3209), .B0(n3211), .B1(n427), .Y(n1834) );
  OAI22XL U2509 ( .A0(n3116), .A1(n3207), .B0(n3206), .B1(n402), .Y(n1859) );
  OAI22XL U2510 ( .A0(n3114), .A1(n3204), .B0(n3206), .B1(n401), .Y(n1860) );
  OAI22XL U2511 ( .A0(n3112), .A1(n3204), .B0(n3206), .B1(n400), .Y(n1861) );
  OAI22XL U2512 ( .A0(n3110), .A1(n3207), .B0(n3206), .B1(n399), .Y(n1862) );
  OAI22XL U2513 ( .A0(n3108), .A1(n3204), .B0(n3206), .B1(n398), .Y(n1863) );
  OAI22XL U2514 ( .A0(n3106), .A1(n3207), .B0(n3206), .B1(n397), .Y(n1864) );
  OAI22XL U2515 ( .A0(n3104), .A1(n3204), .B0(n3206), .B1(n396), .Y(n1865) );
  OAI22XL U2516 ( .A0(n3102), .A1(n3204), .B0(n3206), .B1(n395), .Y(n1866) );
  OAI22XL U2517 ( .A0(n3116), .A1(n3200), .B0(n3201), .B1(n370), .Y(n1891) );
  OAI22XL U2518 ( .A0(n3114), .A1(n3200), .B0(n3202), .B1(n369), .Y(n1892) );
  OAI22XL U2519 ( .A0(n3112), .A1(n3200), .B0(n3201), .B1(n368), .Y(n1893) );
  OAI22XL U2520 ( .A0(n3110), .A1(n104), .B0(n3202), .B1(n367), .Y(n1894) );
  OAI22XL U2521 ( .A0(n3108), .A1(n3200), .B0(n3201), .B1(n366), .Y(n1895) );
  OAI22XL U2522 ( .A0(n3106), .A1(n3203), .B0(n3202), .B1(n365), .Y(n1896) );
  OAI22XL U2523 ( .A0(n3104), .A1(n3203), .B0(n3201), .B1(n364), .Y(n1897) );
  OAI22XL U2524 ( .A0(n3102), .A1(n3200), .B0(n3202), .B1(n363), .Y(n1898) );
  OAI22XL U2525 ( .A0(n3116), .A1(n3199), .B0(n3197), .B1(n338), .Y(n1923) );
  OAI22XL U2526 ( .A0(n3114), .A1(n3196), .B0(n3198), .B1(n337), .Y(n1924) );
  OAI22XL U2527 ( .A0(n3112), .A1(n3199), .B0(n3197), .B1(n336), .Y(n1925) );
  OAI22XL U2528 ( .A0(n3110), .A1(n3196), .B0(n3198), .B1(n335), .Y(n1926) );
  OAI22XL U2529 ( .A0(n3108), .A1(n3196), .B0(n3197), .B1(n334), .Y(n1927) );
  OAI22XL U2530 ( .A0(n3106), .A1(n3196), .B0(n3198), .B1(n333), .Y(n1928) );
  OAI22XL U2531 ( .A0(n3104), .A1(n3199), .B0(n3197), .B1(n332), .Y(n1929) );
  OAI22XL U2532 ( .A0(n3102), .A1(n3199), .B0(n3198), .B1(n331), .Y(n1930) );
  OAI22XL U2533 ( .A0(n3116), .A1(n3192), .B0(n3193), .B1(n306), .Y(n1955) );
  OAI22XL U2534 ( .A0(n3114), .A1(n3192), .B0(n3194), .B1(n305), .Y(n1956) );
  OAI22XL U2535 ( .A0(n3112), .A1(n3192), .B0(n3193), .B1(n304), .Y(n1957) );
  OAI22XL U2536 ( .A0(n3110), .A1(n110), .B0(n3194), .B1(n303), .Y(n1958) );
  OAI22XL U2537 ( .A0(n3108), .A1(n3192), .B0(n3193), .B1(n302), .Y(n1959) );
  OAI22XL U2538 ( .A0(n3106), .A1(n3195), .B0(n3194), .B1(n301), .Y(n1960) );
  OAI22XL U2539 ( .A0(n3104), .A1(n3195), .B0(n3193), .B1(n300), .Y(n1961) );
  OAI22XL U2540 ( .A0(n3102), .A1(n3192), .B0(n3194), .B1(n299), .Y(n1962) );
  OAI22XL U2541 ( .A0(n3116), .A1(n3191), .B0(n3189), .B1(n274), .Y(n1987) );
  OAI22XL U2542 ( .A0(n3114), .A1(n3188), .B0(n3190), .B1(n273), .Y(n1988) );
  OAI22XL U2543 ( .A0(n3112), .A1(n3191), .B0(n3189), .B1(n272), .Y(n1989) );
  OAI22XL U2544 ( .A0(n3110), .A1(n3188), .B0(n3190), .B1(n271), .Y(n1990) );
  OAI22XL U2545 ( .A0(n3108), .A1(n3188), .B0(n3189), .B1(n270), .Y(n1991) );
  OAI22XL U2546 ( .A0(n3106), .A1(n3188), .B0(n3190), .B1(n269), .Y(n1992) );
  OAI22XL U2547 ( .A0(n3104), .A1(n3191), .B0(n3189), .B1(n268), .Y(n1993) );
  OAI22XL U2548 ( .A0(n3102), .A1(n3191), .B0(n3190), .B1(n267), .Y(n1994) );
  OAI22XL U2549 ( .A0(n3116), .A1(n3184), .B0(n3185), .B1(n242), .Y(n2019) );
  OAI22XL U2550 ( .A0(n3114), .A1(n3184), .B0(n3186), .B1(n241), .Y(n2020) );
  OAI22XL U2551 ( .A0(n3112), .A1(n3184), .B0(n3185), .B1(n240), .Y(n2021) );
  OAI22XL U2552 ( .A0(n3110), .A1(n115), .B0(n3186), .B1(n239), .Y(n2022) );
  OAI22XL U2553 ( .A0(n3108), .A1(n3184), .B0(n3185), .B1(n238), .Y(n2023) );
  OAI22XL U2554 ( .A0(n3106), .A1(n3187), .B0(n3186), .B1(n237), .Y(n2024) );
  OAI22XL U2555 ( .A0(n3104), .A1(n3187), .B0(n3185), .B1(n236), .Y(n2025) );
  OAI22XL U2556 ( .A0(n3102), .A1(n3184), .B0(n3186), .B1(n235), .Y(n2026) );
  OAI22XL U2557 ( .A0(n3116), .A1(n3183), .B0(n3181), .B1(n210), .Y(n2051) );
  OAI22XL U2558 ( .A0(n3114), .A1(n3180), .B0(n3182), .B1(n209), .Y(n2052) );
  OAI22XL U2559 ( .A0(n3112), .A1(n3183), .B0(n3181), .B1(n208), .Y(n2053) );
  OAI22XL U2560 ( .A0(n3110), .A1(n3180), .B0(n3182), .B1(n207), .Y(n2054) );
  OAI22XL U2561 ( .A0(n3108), .A1(n3180), .B0(n3181), .B1(n206), .Y(n2055) );
  OAI22XL U2562 ( .A0(n3106), .A1(n3180), .B0(n3182), .B1(n205), .Y(n2056) );
  OAI22XL U2563 ( .A0(n3104), .A1(n3183), .B0(n3181), .B1(n204), .Y(n2057) );
  OAI22XL U2564 ( .A0(n3102), .A1(n3183), .B0(n3182), .B1(n203), .Y(n2058) );
  OAI22XL U2565 ( .A0(n3116), .A1(n3176), .B0(n3177), .B1(n178), .Y(n2083) );
  OAI22XL U2566 ( .A0(n3114), .A1(n3176), .B0(n3178), .B1(n177), .Y(n2084) );
  OAI22XL U2567 ( .A0(n3112), .A1(n3176), .B0(n3177), .B1(n176), .Y(n2085) );
  OAI22XL U2568 ( .A0(n3110), .A1(n120), .B0(n3178), .B1(n175), .Y(n2086) );
  OAI22XL U2569 ( .A0(n3108), .A1(n3176), .B0(n3177), .B1(n174), .Y(n2087) );
  OAI22XL U2570 ( .A0(n3106), .A1(n3179), .B0(n3178), .B1(n173), .Y(n2088) );
  OAI22XL U2571 ( .A0(n3104), .A1(n3179), .B0(n3177), .B1(n172), .Y(n2089) );
  OAI22XL U2572 ( .A0(n3102), .A1(n3176), .B0(n3178), .B1(n171), .Y(n2090) );
  OAI22XL U2573 ( .A0(n3116), .A1(n3175), .B0(n3173), .B1(n146), .Y(n2115) );
  OAI22XL U2574 ( .A0(n3114), .A1(n3172), .B0(n3174), .B1(n145), .Y(n2116) );
  OAI22XL U2575 ( .A0(n3112), .A1(n3175), .B0(n3173), .B1(n144), .Y(n2117) );
  OAI22XL U2576 ( .A0(n3110), .A1(n3172), .B0(n3174), .B1(n143), .Y(n2118) );
  OAI22XL U2577 ( .A0(n3108), .A1(n3172), .B0(n3173), .B1(n142), .Y(n2119) );
  OAI22XL U2578 ( .A0(n3106), .A1(n3172), .B0(n3174), .B1(n141), .Y(n2120) );
  OAI22XL U2579 ( .A0(n3104), .A1(n3175), .B0(n3173), .B1(n140), .Y(n2121) );
  OAI22XL U2580 ( .A0(n3102), .A1(n3175), .B0(n3174), .B1(n139), .Y(n2122) );
  NOR2BX1 U2581 ( .AN(n103), .B(WriteReg[3]), .Y(n100) );
  AND2X2 U2582 ( .A(WriteReg[4]), .B(RegWrite), .Y(n103) );
endmodule


module aluCtrl ( opcode, funct, ALUOp, ctrl );
  input [5:0] opcode;
  input [5:0] funct;
  input [1:0] ALUOp;
  output [3:0] ctrl;
  wire   n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n1, n2, n3, n4, n5, n6, n7, n8, n9, n41;

  OAI211X2 U9 ( .A0(n41), .A1(n23), .B0(n24), .C0(n25), .Y(ctrl[1]) );
  OAI211X2 U14 ( .A0(n1), .A1(n33), .B0(n2), .C0(n11), .Y(ctrl[0]) );
  CLKINVX1 U2 ( .A(n29), .Y(n6) );
  OA21XL U3 ( .A0(n41), .A1(n32), .B0(n25), .Y(n11) );
  OAI22XL U4 ( .A0(n6), .A1(n38), .B0(n7), .B1(n29), .Y(n14) );
  OAI21XL U5 ( .A0(n6), .A1(n30), .B0(n38), .Y(n27) );
  CLKINVX1 U6 ( .A(n30), .Y(n7) );
  CLKINVX1 U7 ( .A(n20), .Y(n8) );
  AO22X1 U8 ( .A0(opcode[5]), .A1(n1), .B0(funct[5]), .B1(n41), .Y(n29) );
  AOI22X1 U10 ( .A0(opcode[4]), .A1(n1), .B0(funct[4]), .B1(n41), .Y(n38) );
  AO22X1 U11 ( .A0(opcode[2]), .A1(n1), .B0(funct[2]), .B1(n41), .Y(n30) );
  AO22X1 U12 ( .A0(opcode[3]), .A1(n1), .B0(funct[3]), .B1(n41), .Y(n16) );
  OAI211X1 U13 ( .A0(n34), .A1(n17), .B0(n35), .C0(n2), .Y(n32) );
  CLKINVX1 U15 ( .A(n15), .Y(n5) );
  CLKINVX1 U16 ( .A(n35), .Y(n4) );
  AOI211X1 U17 ( .A0(n8), .A1(n12), .B0(n39), .C0(n3), .Y(n33) );
  AO22X1 U18 ( .A0(n9), .A1(n5), .B0(n20), .B1(n22), .Y(n39) );
  OAI31XL U19 ( .A0(n26), .A1(n16), .A2(n27), .B0(n41), .Y(n24) );
  AND3X2 U20 ( .A(n31), .B(n32), .C(n30), .Y(n23) );
  OAI32X1 U21 ( .A0(n12), .A1(n8), .A2(n6), .B0(n28), .B1(n29), .Y(n26) );
  OAI211X1 U22 ( .A0(n1), .A1(n18), .B0(n19), .C0(n11), .Y(ctrl[2]) );
  NAND3X1 U23 ( .A(n4), .B(n20), .C(n7), .Y(n19) );
  AOI211X1 U24 ( .A0(n8), .A1(n5), .B0(n3), .C0(n21), .Y(n18) );
  NOR3X1 U25 ( .A(n22), .B(n8), .C(n6), .Y(n21) );
  CLKINVX1 U26 ( .A(n12), .Y(n9) );
  NAND2X1 U27 ( .A(n6), .B(n38), .Y(n15) );
  NAND2X1 U28 ( .A(n4), .B(n20), .Y(n31) );
  NAND3X1 U29 ( .A(n9), .B(n16), .C(n5), .Y(n35) );
  CLKINVX1 U30 ( .A(n36), .Y(n2) );
  OAI31XL U31 ( .A0(n37), .A1(n34), .A2(n20), .B0(n31), .Y(n36) );
  NAND3X1 U32 ( .A(n16), .B(n30), .C(n6), .Y(n37) );
  INVX3 U33 ( .A(n1), .Y(n41) );
  OAI21X1 U34 ( .A0(n1), .A1(n10), .B0(n11), .Y(ctrl[3]) );
  AOI211X1 U35 ( .A0(n7), .A1(n12), .B0(n13), .C0(n14), .Y(n10) );
  OAI2BB2XL U36 ( .B0(n8), .B1(n15), .A0N(n16), .A1N(n17), .Y(n13) );
  CLKINVX1 U37 ( .A(n40), .Y(n3) );
  AOI211X1 U38 ( .A0(n12), .A1(n27), .B0(n14), .C0(n16), .Y(n40) );
  NOR2X1 U39 ( .A(n12), .B(n7), .Y(n22) );
  NAND2X1 U40 ( .A(n38), .B(n12), .Y(n34) );
  NAND3X1 U41 ( .A(n29), .B(n20), .C(n7), .Y(n17) );
  AOI2BB1X1 U42 ( .A0N(n20), .A1N(n9), .B0(n30), .Y(n28) );
  AO22X2 U43 ( .A0(opcode[0]), .A1(n1), .B0(funct[0]), .B1(n41), .Y(n12) );
  CLKBUFX3 U44 ( .A(ALUOp[0]), .Y(n1) );
  AO22X2 U45 ( .A0(opcode[1]), .A1(n1), .B0(funct[1]), .B1(n41), .Y(n20) );
  XOR2X1 U46 ( .A(n1), .B(ALUOp[1]), .Y(n25) );
endmodule


module alu_DW_rightsh_0 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488;

  NAND4X1 U256 ( .A(n478), .B(n479), .C(n480), .D(n481), .Y(n323) );
  MXI3X1 U257 ( .A(n392), .B(n393), .C(n351), .S0(n328), .S1(n325), .Y(n324)
         );
  CLKBUFX3 U258 ( .A(SH[2]), .Y(n325) );
  CLKINVX1 U259 ( .A(SH[1]), .Y(n356) );
  CLKINVX1 U260 ( .A(SH[3]), .Y(n353) );
  INVX3 U261 ( .A(n335), .Y(n332) );
  INVX3 U262 ( .A(n335), .Y(n333) );
  CLKINVX1 U263 ( .A(n413), .Y(n342) );
  CLKINVX1 U264 ( .A(n415), .Y(n343) );
  CLKINVX1 U265 ( .A(n417), .Y(n344) );
  CLKINVX1 U266 ( .A(n364), .Y(n348) );
  CLKINVX1 U267 ( .A(n427), .Y(n345) );
  CLKINVX1 U268 ( .A(n429), .Y(n346) );
  CLKINVX1 U269 ( .A(n360), .Y(n347) );
  CLKINVX1 U270 ( .A(n407), .Y(n340) );
  CLKBUFX3 U271 ( .A(n323), .Y(n331) );
  CLKBUFX3 U272 ( .A(n335), .Y(n334) );
  CLKINVX1 U273 ( .A(n382), .Y(n349) );
  INVX4 U274 ( .A(n325), .Y(n355) );
  CLKBUFX3 U275 ( .A(n356), .Y(n328) );
  CLKBUFX3 U276 ( .A(n356), .Y(n329) );
  CLKBUFX3 U277 ( .A(n353), .Y(n326) );
  CLKBUFX3 U278 ( .A(n353), .Y(n327) );
  CLKBUFX3 U279 ( .A(n323), .Y(n330) );
  CLKINVX1 U280 ( .A(SH[0]), .Y(n335) );
  CLKBUFX3 U281 ( .A(SH[4]), .Y(n337) );
  CLKBUFX3 U282 ( .A(SH[4]), .Y(n336) );
  CLKBUFX3 U283 ( .A(SH[5]), .Y(n339) );
  CLKINVX1 U284 ( .A(n405), .Y(n352) );
  CLKINVX1 U285 ( .A(n369), .Y(n351) );
  CLKINVX1 U286 ( .A(n403), .Y(n354) );
  CLKINVX1 U287 ( .A(n385), .Y(n341) );
  CLKINVX1 U288 ( .A(n388), .Y(n350) );
  CLKBUFX3 U289 ( .A(SH[5]), .Y(n338) );
  NOR3X1 U290 ( .A(n357), .B(n339), .C(n331), .Y(B[9]) );
  MX3XL U291 ( .A(n347), .B(n358), .C(n359), .S0(n326), .S1(n336), .Y(n357) );
  NOR3X1 U292 ( .A(n361), .B(n338), .C(n331), .Y(B[8]) );
  MX3XL U293 ( .A(n348), .B(n362), .C(n363), .S0(n326), .S1(n336), .Y(n361) );
  NOR3X1 U294 ( .A(n365), .B(n338), .C(n331), .Y(B[7]) );
  CLKMX2X2 U295 ( .A(n366), .B(n367), .S0(n336), .Y(n365) );
  MX3XL U296 ( .A(n368), .B(n369), .C(n370), .S0(n355), .S1(SH[3]), .Y(n366)
         );
  NOR3X1 U297 ( .A(n371), .B(n338), .C(n331), .Y(B[6]) );
  CLKMX2X2 U298 ( .A(n372), .B(n373), .S0(n336), .Y(n371) );
  MX3XL U299 ( .A(n374), .B(n375), .C(n376), .S0(n355), .S1(SH[3]), .Y(n372)
         );
  NOR3X1 U300 ( .A(n377), .B(n338), .C(n331), .Y(B[5]) );
  MX3XL U301 ( .A(n378), .B(n379), .C(n380), .S0(n327), .S1(n337), .Y(n377) );
  MXI2X1 U302 ( .A(n349), .B(n381), .S0(n355), .Y(n379) );
  NOR3X1 U303 ( .A(n383), .B(n338), .C(n331), .Y(B[4]) );
  MXI2X1 U304 ( .A(n384), .B(n341), .S0(n336), .Y(n383) );
  MX3XL U305 ( .A(n350), .B(n386), .C(n387), .S0(n355), .S1(SH[3]), .Y(n384)
         );
  NOR3X1 U306 ( .A(n389), .B(n338), .C(n331), .Y(B[3]) );
  MX3XL U307 ( .A(n390), .B(n324), .C(n391), .S0(n327), .S1(n337), .Y(n389) );
  MXI2X1 U308 ( .A(n394), .B(n395), .S0(n328), .Y(n369) );
  NOR4X1 U309 ( .A(SH[5]), .B(n337), .C(n330), .D(n396), .Y(B[31]) );
  NOR4X1 U310 ( .A(SH[5]), .B(n337), .C(n330), .D(n397), .Y(B[30]) );
  NOR3X1 U311 ( .A(n398), .B(n339), .C(n331), .Y(B[2]) );
  MX3XL U312 ( .A(n399), .B(n400), .C(n401), .S0(n326), .S1(n337), .Y(n398) );
  MX3XL U313 ( .A(n402), .B(n403), .C(n375), .S0(n329), .S1(n325), .Y(n400) );
  MXI2X1 U314 ( .A(n404), .B(n352), .S0(n328), .Y(n375) );
  NOR4X1 U315 ( .A(n338), .B(n337), .C(n330), .D(n406), .Y(B[29]) );
  NOR4X1 U316 ( .A(n339), .B(n337), .C(n330), .D(n407), .Y(B[28]) );
  NOR4X1 U317 ( .A(n339), .B(n337), .C(n330), .D(n408), .Y(B[27]) );
  NOR4X1 U318 ( .A(SH[5]), .B(n337), .C(n330), .D(n409), .Y(B[26]) );
  NOR4X1 U319 ( .A(n339), .B(n337), .C(n330), .D(n359), .Y(B[25]) );
  NAND2X1 U320 ( .A(n410), .B(n327), .Y(n359) );
  NOR4X1 U321 ( .A(SH[5]), .B(n337), .C(n330), .D(n363), .Y(B[24]) );
  NAND2X1 U322 ( .A(n411), .B(n327), .Y(n363) );
  NOR4X1 U323 ( .A(n339), .B(n337), .C(n367), .D(n331), .Y(B[23]) );
  MXI2X1 U324 ( .A(n412), .B(n413), .S0(n326), .Y(n367) );
  NOR4X1 U325 ( .A(SH[5]), .B(n337), .C(n373), .D(n331), .Y(B[22]) );
  MXI2X1 U326 ( .A(n414), .B(n415), .S0(n326), .Y(n373) );
  NOR4X1 U327 ( .A(n339), .B(n337), .C(n380), .D(n331), .Y(B[21]) );
  MXI2X1 U328 ( .A(n416), .B(n417), .S0(n326), .Y(n380) );
  NOR4X1 U329 ( .A(n339), .B(n337), .C(n385), .D(n330), .Y(B[20]) );
  MXI2X1 U330 ( .A(n418), .B(n419), .S0(n326), .Y(n385) );
  NOR3X1 U331 ( .A(n420), .B(n339), .C(n331), .Y(B[1]) );
  MX3XL U332 ( .A(n358), .B(n421), .C(n422), .S0(n326), .S1(n336), .Y(n420) );
  MXI2X1 U333 ( .A(n381), .B(n423), .S0(n355), .Y(n421) );
  MX3XL U334 ( .A(A[2]), .B(A[1]), .C(n393), .S0(n334), .S1(SH[1]), .Y(n423)
         );
  CLKMX2X2 U335 ( .A(A[3]), .B(A[4]), .S0(n332), .Y(n393) );
  CLKMX2X2 U336 ( .A(n392), .B(n395), .S0(SH[1]), .Y(n381) );
  CLKMX2X2 U337 ( .A(A[7]), .B(A[8]), .S0(n332), .Y(n395) );
  CLKMX2X2 U338 ( .A(A[5]), .B(A[6]), .S0(n332), .Y(n392) );
  CLKMX2X2 U339 ( .A(n382), .B(n424), .S0(n325), .Y(n358) );
  MXI2X1 U340 ( .A(n425), .B(n394), .S0(n328), .Y(n382) );
  CLKMX2X2 U341 ( .A(A[9]), .B(A[10]), .S0(n332), .Y(n394) );
  NOR4X1 U342 ( .A(n339), .B(n337), .C(n391), .D(n330), .Y(B[19]) );
  MXI2X1 U343 ( .A(n426), .B(n427), .S0(n326), .Y(n391) );
  NOR4X1 U344 ( .A(n339), .B(n337), .C(n401), .D(n330), .Y(B[18]) );
  MXI2X1 U345 ( .A(n428), .B(n429), .S0(n326), .Y(n401) );
  NOR4X1 U346 ( .A(SH[5]), .B(n337), .C(n422), .D(n330), .Y(B[17]) );
  MXI2X1 U347 ( .A(n410), .B(n360), .S0(n326), .Y(n422) );
  MXI2X1 U348 ( .A(n430), .B(n431), .S0(n355), .Y(n360) );
  MXI2X1 U349 ( .A(n432), .B(n433), .S0(n355), .Y(n410) );
  NOR4X1 U350 ( .A(SH[5]), .B(SH[4]), .C(n434), .D(n330), .Y(B[16]) );
  NOR3X1 U351 ( .A(n435), .B(n339), .C(n330), .Y(B[15]) );
  MX3XL U352 ( .A(n342), .B(n370), .C(n396), .S0(n327), .S1(n336), .Y(n435) );
  NAND2X1 U353 ( .A(n412), .B(n327), .Y(n396) );
  NOR2X1 U354 ( .A(n436), .B(n325), .Y(n412) );
  CLKMX2X2 U355 ( .A(n437), .B(n438), .S0(n325), .Y(n370) );
  MXI2X1 U356 ( .A(n439), .B(n440), .S0(n355), .Y(n413) );
  NOR3X1 U357 ( .A(n441), .B(n339), .C(n323), .Y(B[14]) );
  MX3XL U358 ( .A(n343), .B(n376), .C(n397), .S0(n327), .S1(n336), .Y(n441) );
  NAND2X1 U359 ( .A(n414), .B(n327), .Y(n397) );
  NOR2X1 U360 ( .A(n442), .B(n325), .Y(n414) );
  CLKMX2X2 U361 ( .A(n443), .B(n444), .S0(n325), .Y(n376) );
  MXI2X1 U362 ( .A(n445), .B(n446), .S0(n355), .Y(n415) );
  NOR3X1 U363 ( .A(n447), .B(n339), .C(n323), .Y(B[13]) );
  MX3XL U364 ( .A(n344), .B(n378), .C(n406), .S0(n327), .S1(n336), .Y(n447) );
  NAND2X1 U365 ( .A(n416), .B(n327), .Y(n406) );
  NOR2X1 U366 ( .A(n432), .B(n325), .Y(n416) );
  MXI2X1 U367 ( .A(n448), .B(n449), .S0(n328), .Y(n432) );
  CLKMX2X2 U368 ( .A(n424), .B(n431), .S0(n325), .Y(n378) );
  MXI2X1 U369 ( .A(n450), .B(n451), .S0(n329), .Y(n431) );
  MXI2X1 U370 ( .A(n452), .B(n453), .S0(n328), .Y(n424) );
  MXI2X1 U371 ( .A(n433), .B(n430), .S0(n355), .Y(n417) );
  MXI2X1 U372 ( .A(n454), .B(n455), .S0(n328), .Y(n430) );
  MXI2X1 U373 ( .A(n456), .B(n457), .S0(n328), .Y(n433) );
  NOR3BXL U374 ( .AN(n458), .B(n338), .C(n323), .Y(B[12]) );
  MX3XL U375 ( .A(n419), .B(n387), .C(n340), .S0(n327), .S1(n336), .Y(n458) );
  NAND2X1 U376 ( .A(n418), .B(n327), .Y(n407) );
  NOR2X1 U377 ( .A(n459), .B(n325), .Y(n418) );
  MXI2X1 U378 ( .A(n460), .B(n461), .S0(n355), .Y(n387) );
  MXI2X1 U379 ( .A(n462), .B(n463), .S0(n355), .Y(n419) );
  NOR3X1 U380 ( .A(n464), .B(n339), .C(n323), .Y(B[11]) );
  MX3XL U381 ( .A(n345), .B(n390), .C(n408), .S0(n327), .S1(n336), .Y(n464) );
  NAND2X1 U382 ( .A(n426), .B(n326), .Y(n408) );
  MXI2X1 U383 ( .A(n436), .B(n439), .S0(n355), .Y(n426) );
  MXI2X1 U384 ( .A(n449), .B(n456), .S0(n328), .Y(n439) );
  CLKMX2X2 U385 ( .A(A[27]), .B(A[28]), .S0(n332), .Y(n456) );
  CLKMX2X2 U386 ( .A(A[29]), .B(A[30]), .S0(n332), .Y(n449) );
  NAND2X1 U387 ( .A(n448), .B(n328), .Y(n436) );
  AND2X1 U388 ( .A(A[31]), .B(n334), .Y(n448) );
  CLKMX2X2 U389 ( .A(n368), .B(n437), .S0(n325), .Y(n390) );
  MXI2X1 U390 ( .A(n451), .B(n452), .S0(n328), .Y(n437) );
  CLKMX2X2 U391 ( .A(A[15]), .B(A[16]), .S0(n332), .Y(n452) );
  CLKMX2X2 U392 ( .A(A[17]), .B(A[18]), .S0(n332), .Y(n451) );
  MXI2X1 U393 ( .A(n453), .B(n425), .S0(n328), .Y(n368) );
  CLKMX2X2 U394 ( .A(A[11]), .B(A[12]), .S0(n332), .Y(n425) );
  CLKMX2X2 U395 ( .A(A[13]), .B(A[14]), .S0(n332), .Y(n453) );
  MXI2X1 U396 ( .A(n440), .B(n438), .S0(n355), .Y(n427) );
  MXI2X1 U397 ( .A(n455), .B(n450), .S0(n328), .Y(n438) );
  CLKMX2X2 U398 ( .A(A[19]), .B(A[20]), .S0(n332), .Y(n450) );
  CLKMX2X2 U399 ( .A(A[21]), .B(A[22]), .S0(n332), .Y(n455) );
  MXI2X1 U400 ( .A(n457), .B(n454), .S0(n328), .Y(n440) );
  CLKMX2X2 U401 ( .A(A[23]), .B(A[24]), .S0(n332), .Y(n454) );
  CLKMX2X2 U402 ( .A(A[25]), .B(A[26]), .S0(n333), .Y(n457) );
  NOR3X1 U403 ( .A(n465), .B(n339), .C(n331), .Y(B[10]) );
  MX3XL U404 ( .A(n346), .B(n399), .C(n409), .S0(n327), .S1(n336), .Y(n465) );
  NAND2X1 U405 ( .A(n428), .B(n327), .Y(n409) );
  MXI2X1 U406 ( .A(n442), .B(n445), .S0(n355), .Y(n428) );
  MXI2X1 U407 ( .A(n466), .B(n467), .S0(n329), .Y(n445) );
  NAND2X1 U408 ( .A(n468), .B(n328), .Y(n442) );
  CLKMX2X2 U409 ( .A(n374), .B(n443), .S0(n325), .Y(n399) );
  MXI2X1 U410 ( .A(n469), .B(n470), .S0(n329), .Y(n443) );
  MXI2X1 U411 ( .A(n471), .B(n472), .S0(n329), .Y(n374) );
  MXI2X1 U412 ( .A(n446), .B(n444), .S0(n355), .Y(n429) );
  MXI2X1 U413 ( .A(n473), .B(n474), .S0(n329), .Y(n444) );
  MXI2X1 U414 ( .A(n475), .B(n476), .S0(n329), .Y(n446) );
  NOR3X1 U415 ( .A(n477), .B(n339), .C(n331), .Y(B[0]) );
  AND4X1 U416 ( .A(n482), .B(n483), .C(n484), .D(n485), .Y(n481) );
  NOR4X1 U417 ( .A(SH[9]), .B(SH[8]), .C(SH[7]), .D(SH[6]), .Y(n485) );
  NOR3X1 U418 ( .A(SH[29]), .B(SH[31]), .C(SH[30]), .Y(n484) );
  NOR3X1 U419 ( .A(SH[26]), .B(SH[28]), .C(SH[27]), .Y(n483) );
  NOR3X1 U420 ( .A(SH[23]), .B(SH[25]), .C(SH[24]), .Y(n482) );
  NOR4X1 U421 ( .A(n486), .B(SH[16]), .C(SH[18]), .D(SH[17]), .Y(n480) );
  OR4X1 U422 ( .A(SH[20]), .B(SH[19]), .C(SH[22]), .D(SH[21]), .Y(n486) );
  NOR3X1 U423 ( .A(SH[13]), .B(SH[15]), .C(SH[14]), .Y(n479) );
  NOR3X1 U424 ( .A(SH[10]), .B(SH[12]), .C(SH[11]), .Y(n478) );
  MX3XL U425 ( .A(n362), .B(n487), .C(n434), .S0(n326), .S1(n336), .Y(n477) );
  MXI2X1 U426 ( .A(n411), .B(n364), .S0(n326), .Y(n434) );
  MXI2X1 U427 ( .A(n463), .B(n460), .S0(n355), .Y(n364) );
  MXI2X1 U428 ( .A(n474), .B(n469), .S0(n329), .Y(n460) );
  CLKMX2X2 U429 ( .A(A[16]), .B(A[17]), .S0(n333), .Y(n469) );
  CLKMX2X2 U430 ( .A(A[18]), .B(A[19]), .S0(n333), .Y(n474) );
  MXI2X1 U431 ( .A(n476), .B(n473), .S0(n329), .Y(n463) );
  CLKMX2X2 U432 ( .A(A[20]), .B(A[21]), .S0(n333), .Y(n473) );
  CLKMX2X2 U433 ( .A(A[22]), .B(A[23]), .S0(n333), .Y(n476) );
  MXI2X1 U434 ( .A(n459), .B(n462), .S0(n355), .Y(n411) );
  MXI2X1 U435 ( .A(n467), .B(n475), .S0(n329), .Y(n462) );
  CLKMX2X2 U436 ( .A(A[24]), .B(A[25]), .S0(n333), .Y(n475) );
  CLKMX2X2 U437 ( .A(A[26]), .B(A[27]), .S0(n333), .Y(n467) );
  MXI2X1 U438 ( .A(n468), .B(n466), .S0(n329), .Y(n459) );
  CLKMX2X2 U439 ( .A(A[28]), .B(A[29]), .S0(n333), .Y(n466) );
  CLKMX2X2 U440 ( .A(A[30]), .B(A[31]), .S0(n333), .Y(n468) );
  MXI2X1 U441 ( .A(n386), .B(n488), .S0(n355), .Y(n487) );
  MX3XL U442 ( .A(A[1]), .B(A[0]), .C(n354), .S0(n334), .S1(SH[1]), .Y(n488)
         );
  MXI2X1 U443 ( .A(A[3]), .B(A[2]), .S0(n334), .Y(n403) );
  MXI2X1 U444 ( .A(n405), .B(n402), .S0(n329), .Y(n386) );
  MXI2X1 U445 ( .A(A[5]), .B(A[4]), .S0(n334), .Y(n402) );
  MXI2X1 U446 ( .A(A[7]), .B(A[6]), .S0(n334), .Y(n405) );
  CLKMX2X2 U447 ( .A(n388), .B(n461), .S0(n325), .Y(n362) );
  MXI2X1 U448 ( .A(n470), .B(n471), .S0(n329), .Y(n461) );
  CLKMX2X2 U449 ( .A(A[12]), .B(A[13]), .S0(n333), .Y(n471) );
  CLKMX2X2 U450 ( .A(A[14]), .B(A[15]), .S0(n333), .Y(n470) );
  MXI2X1 U451 ( .A(n472), .B(n404), .S0(n328), .Y(n388) );
  CLKMX2X2 U452 ( .A(A[8]), .B(A[9]), .S0(n333), .Y(n404) );
  CLKMX2X2 U453 ( .A(A[10]), .B(A[11]), .S0(n333), .Y(n472) );
endmodule


module alu_DW_rightsh_1 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487;

  NAND4X1 U256 ( .A(n477), .B(n478), .C(n479), .D(n480), .Y(n323) );
  MXI3X1 U257 ( .A(n391), .B(n392), .C(n353), .S0(n337), .S1(n333), .Y(n324)
         );
  CLKINVX1 U258 ( .A(n384), .Y(n343) );
  CLKINVX1 U259 ( .A(n412), .Y(n344) );
  CLKINVX1 U260 ( .A(n414), .Y(n345) );
  CLKINVX1 U261 ( .A(n416), .Y(n346) );
  CLKINVX1 U262 ( .A(n426), .Y(n347) );
  CLKINVX1 U263 ( .A(n428), .Y(n348) );
  CLKINVX1 U264 ( .A(n359), .Y(n349) );
  CLKINVX1 U265 ( .A(n363), .Y(n350) );
  CLKINVX1 U266 ( .A(n406), .Y(n342) );
  CLKINVX1 U267 ( .A(n381), .Y(n351) );
  INVX3 U268 ( .A(n341), .Y(n338) );
  INVX3 U269 ( .A(n341), .Y(n339) );
  INVX3 U270 ( .A(n333), .Y(n334) );
  CLKINVX1 U271 ( .A(SH[2]), .Y(n335) );
  CLKINVX1 U272 ( .A(n404), .Y(n354) );
  CLKINVX1 U273 ( .A(n387), .Y(n352) );
  CLKINVX1 U274 ( .A(n368), .Y(n353) );
  CLKBUFX3 U275 ( .A(n323), .Y(n326) );
  INVX3 U276 ( .A(SH[1]), .Y(n336) );
  INVX3 U277 ( .A(SH[1]), .Y(n337) );
  CLKBUFX3 U278 ( .A(n341), .Y(n340) );
  CLKBUFX3 U279 ( .A(SH[4]), .Y(n330) );
  CLKBUFX3 U280 ( .A(SH[4]), .Y(n329) );
  CLKBUFX3 U281 ( .A(SH[5]), .Y(n328) );
  CLKBUFX3 U282 ( .A(SH[5]), .Y(n327) );
  INVX3 U283 ( .A(SH[3]), .Y(n331) );
  INVX3 U284 ( .A(SH[3]), .Y(n332) );
  CLKINVX1 U285 ( .A(n402), .Y(n355) );
  CLKBUFX3 U286 ( .A(n323), .Y(n325) );
  CLKBUFX3 U287 ( .A(SH[2]), .Y(n333) );
  CLKINVX1 U288 ( .A(SH[0]), .Y(n341) );
  NOR3X1 U289 ( .A(n356), .B(n328), .C(n326), .Y(B[9]) );
  MX3XL U290 ( .A(n349), .B(n357), .C(n358), .S0(n331), .S1(n329), .Y(n356) );
  NOR3X1 U291 ( .A(n360), .B(SH[5]), .C(n326), .Y(B[8]) );
  MX3XL U292 ( .A(n350), .B(n361), .C(n362), .S0(n332), .S1(n329), .Y(n360) );
  NOR3X1 U293 ( .A(n364), .B(SH[5]), .C(n326), .Y(B[7]) );
  CLKMX2X2 U294 ( .A(n365), .B(n366), .S0(n329), .Y(n364) );
  MX3XL U295 ( .A(n367), .B(n368), .C(n369), .S0(n335), .S1(SH[3]), .Y(n365)
         );
  NOR3X1 U296 ( .A(n370), .B(SH[5]), .C(n326), .Y(B[6]) );
  CLKMX2X2 U297 ( .A(n371), .B(n372), .S0(n329), .Y(n370) );
  MX3XL U298 ( .A(n373), .B(n374), .C(n375), .S0(n335), .S1(SH[3]), .Y(n371)
         );
  NOR3X1 U299 ( .A(n376), .B(SH[5]), .C(n326), .Y(B[5]) );
  MX3XL U300 ( .A(n377), .B(n378), .C(n379), .S0(n332), .S1(n330), .Y(n376) );
  MXI2X1 U301 ( .A(n351), .B(n380), .S0(n335), .Y(n378) );
  NOR3X1 U302 ( .A(n382), .B(SH[5]), .C(n326), .Y(B[4]) );
  MXI2X1 U303 ( .A(n383), .B(n343), .S0(n329), .Y(n382) );
  MX3XL U304 ( .A(n352), .B(n385), .C(n386), .S0(n335), .S1(SH[3]), .Y(n383)
         );
  NOR3X1 U305 ( .A(n388), .B(n327), .C(n326), .Y(B[3]) );
  MX3XL U306 ( .A(n389), .B(n324), .C(n390), .S0(n332), .S1(n330), .Y(n388) );
  MXI2X1 U307 ( .A(n393), .B(n394), .S0(n337), .Y(n368) );
  NOR4X1 U308 ( .A(n327), .B(n330), .C(n325), .D(n395), .Y(B[31]) );
  NOR4X1 U309 ( .A(n327), .B(n330), .C(n325), .D(n396), .Y(B[30]) );
  NOR3X1 U310 ( .A(n397), .B(n328), .C(n326), .Y(B[2]) );
  MX3XL U311 ( .A(n398), .B(n399), .C(n400), .S0(n332), .S1(n330), .Y(n397) );
  MX3XL U312 ( .A(n401), .B(n402), .C(n374), .S0(n337), .S1(SH[2]), .Y(n399)
         );
  MXI2X1 U313 ( .A(n403), .B(n354), .S0(n337), .Y(n374) );
  NOR4X1 U314 ( .A(n327), .B(n330), .C(n325), .D(n405), .Y(B[29]) );
  NOR4X1 U315 ( .A(n327), .B(n330), .C(n325), .D(n406), .Y(B[28]) );
  NOR4X1 U316 ( .A(n327), .B(n330), .C(n325), .D(n407), .Y(B[27]) );
  NOR4X1 U317 ( .A(n327), .B(n330), .C(n325), .D(n408), .Y(B[26]) );
  NOR4X1 U318 ( .A(n327), .B(n330), .C(n325), .D(n358), .Y(B[25]) );
  NAND2X1 U319 ( .A(n409), .B(n332), .Y(n358) );
  NOR4X1 U320 ( .A(n327), .B(n330), .C(n325), .D(n362), .Y(B[24]) );
  NAND2X1 U321 ( .A(n410), .B(n332), .Y(n362) );
  NOR4X1 U322 ( .A(n328), .B(n330), .C(n366), .D(n326), .Y(B[23]) );
  MXI2X1 U323 ( .A(n411), .B(n412), .S0(n331), .Y(n366) );
  NOR4X1 U324 ( .A(n327), .B(n330), .C(n372), .D(n326), .Y(B[22]) );
  MXI2X1 U325 ( .A(n413), .B(n414), .S0(n331), .Y(n372) );
  NOR4X1 U326 ( .A(n328), .B(n330), .C(n379), .D(n326), .Y(B[21]) );
  MXI2X1 U327 ( .A(n415), .B(n416), .S0(n331), .Y(n379) );
  NOR4X1 U328 ( .A(n328), .B(n330), .C(n384), .D(n325), .Y(B[20]) );
  MXI2X1 U329 ( .A(n417), .B(n418), .S0(n331), .Y(n384) );
  NOR3X1 U330 ( .A(n419), .B(n328), .C(n326), .Y(B[1]) );
  MX3XL U331 ( .A(n357), .B(n420), .C(n421), .S0(n332), .S1(n329), .Y(n419) );
  MXI2X1 U332 ( .A(n380), .B(n422), .S0(n335), .Y(n420) );
  MX3XL U333 ( .A(A[2]), .B(A[1]), .C(n392), .S0(n340), .S1(SH[1]), .Y(n422)
         );
  CLKMX2X2 U334 ( .A(A[3]), .B(A[4]), .S0(n338), .Y(n392) );
  CLKMX2X2 U335 ( .A(n391), .B(n394), .S0(SH[1]), .Y(n380) );
  CLKMX2X2 U336 ( .A(A[7]), .B(A[8]), .S0(n338), .Y(n394) );
  CLKMX2X2 U337 ( .A(A[5]), .B(A[6]), .S0(n338), .Y(n391) );
  CLKMX2X2 U338 ( .A(n381), .B(n423), .S0(n333), .Y(n357) );
  MXI2X1 U339 ( .A(n424), .B(n393), .S0(n337), .Y(n381) );
  CLKMX2X2 U340 ( .A(A[9]), .B(A[10]), .S0(n338), .Y(n393) );
  NOR4X1 U341 ( .A(n327), .B(n330), .C(n390), .D(n325), .Y(B[19]) );
  MXI2X1 U342 ( .A(n425), .B(n426), .S0(n331), .Y(n390) );
  NOR4X1 U343 ( .A(n328), .B(n330), .C(n400), .D(n325), .Y(B[18]) );
  MXI2X1 U344 ( .A(n427), .B(n428), .S0(n331), .Y(n400) );
  NOR4X1 U345 ( .A(n327), .B(n330), .C(n421), .D(n325), .Y(B[17]) );
  MXI2X1 U346 ( .A(n409), .B(n359), .S0(n331), .Y(n421) );
  MXI2X1 U347 ( .A(n429), .B(n430), .S0(n335), .Y(n359) );
  MXI2X1 U348 ( .A(n431), .B(n432), .S0(n334), .Y(n409) );
  NOR4X1 U349 ( .A(n327), .B(SH[4]), .C(n433), .D(n325), .Y(B[16]) );
  NOR3X1 U350 ( .A(n434), .B(n328), .C(n325), .Y(B[15]) );
  MX3XL U351 ( .A(n344), .B(n369), .C(n395), .S0(n331), .S1(n329), .Y(n434) );
  NAND2X1 U352 ( .A(n411), .B(n332), .Y(n395) );
  NOR2X1 U353 ( .A(n435), .B(SH[2]), .Y(n411) );
  CLKMX2X2 U354 ( .A(n436), .B(n437), .S0(SH[2]), .Y(n369) );
  MXI2X1 U355 ( .A(n438), .B(n439), .S0(n334), .Y(n412) );
  NOR3X1 U356 ( .A(n440), .B(n328), .C(n323), .Y(B[14]) );
  MX3XL U357 ( .A(n345), .B(n375), .C(n396), .S0(n332), .S1(n329), .Y(n440) );
  NAND2X1 U358 ( .A(n413), .B(n332), .Y(n396) );
  NOR2X1 U359 ( .A(n441), .B(SH[2]), .Y(n413) );
  CLKMX2X2 U360 ( .A(n442), .B(n443), .S0(SH[2]), .Y(n375) );
  MXI2X1 U361 ( .A(n444), .B(n445), .S0(n334), .Y(n414) );
  NOR3X1 U362 ( .A(n446), .B(n328), .C(n323), .Y(B[13]) );
  MX3XL U363 ( .A(n346), .B(n377), .C(n405), .S0(n331), .S1(n329), .Y(n446) );
  NAND2X1 U364 ( .A(n415), .B(n332), .Y(n405) );
  NOR2X1 U365 ( .A(n431), .B(SH[2]), .Y(n415) );
  MXI2X1 U366 ( .A(n447), .B(n448), .S0(n337), .Y(n431) );
  CLKMX2X2 U367 ( .A(n423), .B(n430), .S0(n333), .Y(n377) );
  MXI2X1 U368 ( .A(n449), .B(n450), .S0(n337), .Y(n430) );
  MXI2X1 U369 ( .A(n451), .B(n452), .S0(n337), .Y(n423) );
  MXI2X1 U370 ( .A(n432), .B(n429), .S0(n334), .Y(n416) );
  MXI2X1 U371 ( .A(n453), .B(n454), .S0(n337), .Y(n429) );
  MXI2X1 U372 ( .A(n455), .B(n456), .S0(n337), .Y(n432) );
  NOR3BXL U373 ( .AN(n457), .B(n327), .C(n323), .Y(B[12]) );
  MX3XL U374 ( .A(n418), .B(n386), .C(n342), .S0(n332), .S1(n329), .Y(n457) );
  NAND2X1 U375 ( .A(n417), .B(n332), .Y(n406) );
  NOR2X1 U376 ( .A(n458), .B(SH[2]), .Y(n417) );
  MXI2X1 U377 ( .A(n459), .B(n460), .S0(n334), .Y(n386) );
  MXI2X1 U378 ( .A(n461), .B(n462), .S0(n334), .Y(n418) );
  NOR3X1 U379 ( .A(n463), .B(n328), .C(n323), .Y(B[11]) );
  MX3XL U380 ( .A(n347), .B(n389), .C(n407), .S0(n331), .S1(n329), .Y(n463) );
  NAND2X1 U381 ( .A(n425), .B(n332), .Y(n407) );
  MXI2X1 U382 ( .A(n435), .B(n438), .S0(n334), .Y(n425) );
  MXI2X1 U383 ( .A(n448), .B(n455), .S0(n337), .Y(n438) );
  CLKMX2X2 U384 ( .A(A[27]), .B(A[28]), .S0(n338), .Y(n455) );
  CLKMX2X2 U385 ( .A(A[29]), .B(A[30]), .S0(n338), .Y(n448) );
  NAND2X1 U386 ( .A(n447), .B(n337), .Y(n435) );
  AND2X1 U387 ( .A(A[31]), .B(n340), .Y(n447) );
  CLKMX2X2 U388 ( .A(n367), .B(n436), .S0(n333), .Y(n389) );
  MXI2X1 U389 ( .A(n450), .B(n451), .S0(n337), .Y(n436) );
  CLKMX2X2 U390 ( .A(A[15]), .B(A[16]), .S0(n338), .Y(n451) );
  CLKMX2X2 U391 ( .A(A[17]), .B(A[18]), .S0(n338), .Y(n450) );
  MXI2X1 U392 ( .A(n452), .B(n424), .S0(n337), .Y(n367) );
  CLKMX2X2 U393 ( .A(A[11]), .B(A[12]), .S0(n338), .Y(n424) );
  CLKMX2X2 U394 ( .A(A[13]), .B(A[14]), .S0(n338), .Y(n452) );
  MXI2X1 U395 ( .A(n439), .B(n437), .S0(n334), .Y(n426) );
  MXI2X1 U396 ( .A(n454), .B(n449), .S0(n336), .Y(n437) );
  CLKMX2X2 U397 ( .A(A[19]), .B(A[20]), .S0(n338), .Y(n449) );
  CLKMX2X2 U398 ( .A(A[21]), .B(A[22]), .S0(n338), .Y(n454) );
  MXI2X1 U399 ( .A(n456), .B(n453), .S0(n336), .Y(n439) );
  CLKMX2X2 U400 ( .A(A[23]), .B(A[24]), .S0(n338), .Y(n453) );
  CLKMX2X2 U401 ( .A(A[25]), .B(A[26]), .S0(n339), .Y(n456) );
  NOR3X1 U402 ( .A(n464), .B(n328), .C(n326), .Y(B[10]) );
  MX3XL U403 ( .A(n348), .B(n398), .C(n408), .S0(n332), .S1(n329), .Y(n464) );
  NAND2X1 U404 ( .A(n427), .B(n331), .Y(n408) );
  MXI2X1 U405 ( .A(n441), .B(n444), .S0(n334), .Y(n427) );
  MXI2X1 U406 ( .A(n465), .B(n466), .S0(n336), .Y(n444) );
  NAND2X1 U407 ( .A(n467), .B(n337), .Y(n441) );
  CLKMX2X2 U408 ( .A(n373), .B(n442), .S0(SH[2]), .Y(n398) );
  MXI2X1 U409 ( .A(n468), .B(n469), .S0(n336), .Y(n442) );
  MXI2X1 U410 ( .A(n470), .B(n471), .S0(n336), .Y(n373) );
  MXI2X1 U411 ( .A(n445), .B(n443), .S0(n334), .Y(n428) );
  MXI2X1 U412 ( .A(n472), .B(n473), .S0(n336), .Y(n443) );
  MXI2X1 U413 ( .A(n474), .B(n475), .S0(n336), .Y(n445) );
  NOR3X1 U414 ( .A(n476), .B(n328), .C(n326), .Y(B[0]) );
  AND4X1 U415 ( .A(n481), .B(n482), .C(n483), .D(n484), .Y(n480) );
  NOR4X1 U416 ( .A(SH[9]), .B(SH[8]), .C(SH[7]), .D(SH[6]), .Y(n484) );
  NOR3X1 U417 ( .A(SH[29]), .B(SH[31]), .C(SH[30]), .Y(n483) );
  NOR3X1 U418 ( .A(SH[26]), .B(SH[28]), .C(SH[27]), .Y(n482) );
  NOR3X1 U419 ( .A(SH[23]), .B(SH[25]), .C(SH[24]), .Y(n481) );
  NOR4X1 U420 ( .A(n485), .B(SH[16]), .C(SH[18]), .D(SH[17]), .Y(n479) );
  OR4X1 U421 ( .A(SH[20]), .B(SH[19]), .C(SH[22]), .D(SH[21]), .Y(n485) );
  NOR3X1 U422 ( .A(SH[13]), .B(SH[15]), .C(SH[14]), .Y(n478) );
  NOR3X1 U423 ( .A(SH[10]), .B(SH[12]), .C(SH[11]), .Y(n477) );
  MX3XL U424 ( .A(n361), .B(n486), .C(n433), .S0(n331), .S1(n329), .Y(n476) );
  MXI2X1 U425 ( .A(n410), .B(n363), .S0(n331), .Y(n433) );
  MXI2X1 U426 ( .A(n462), .B(n459), .S0(n334), .Y(n363) );
  MXI2X1 U427 ( .A(n473), .B(n468), .S0(n336), .Y(n459) );
  CLKMX2X2 U428 ( .A(A[16]), .B(A[17]), .S0(n339), .Y(n468) );
  CLKMX2X2 U429 ( .A(A[18]), .B(A[19]), .S0(n339), .Y(n473) );
  MXI2X1 U430 ( .A(n475), .B(n472), .S0(n336), .Y(n462) );
  CLKMX2X2 U431 ( .A(A[20]), .B(A[21]), .S0(n339), .Y(n472) );
  CLKMX2X2 U432 ( .A(A[22]), .B(A[23]), .S0(n339), .Y(n475) );
  MXI2X1 U433 ( .A(n458), .B(n461), .S0(n334), .Y(n410) );
  MXI2X1 U434 ( .A(n466), .B(n474), .S0(n336), .Y(n461) );
  CLKMX2X2 U435 ( .A(A[24]), .B(A[25]), .S0(n339), .Y(n474) );
  CLKMX2X2 U436 ( .A(A[26]), .B(A[27]), .S0(n339), .Y(n466) );
  MXI2X1 U437 ( .A(n467), .B(n465), .S0(n336), .Y(n458) );
  CLKMX2X2 U438 ( .A(A[28]), .B(A[29]), .S0(n339), .Y(n465) );
  CLKMX2X2 U439 ( .A(A[30]), .B(A[31]), .S0(n339), .Y(n467) );
  MXI2X1 U440 ( .A(n385), .B(n487), .S0(n334), .Y(n486) );
  MX3XL U441 ( .A(A[1]), .B(A[0]), .C(n355), .S0(n340), .S1(SH[1]), .Y(n487)
         );
  MXI2X1 U442 ( .A(A[3]), .B(A[2]), .S0(n340), .Y(n402) );
  MXI2X1 U443 ( .A(n404), .B(n401), .S0(n336), .Y(n385) );
  MXI2X1 U444 ( .A(A[5]), .B(A[4]), .S0(n340), .Y(n401) );
  MXI2X1 U445 ( .A(A[7]), .B(A[6]), .S0(n340), .Y(n404) );
  CLKMX2X2 U446 ( .A(n387), .B(n460), .S0(n333), .Y(n361) );
  MXI2X1 U447 ( .A(n469), .B(n470), .S0(n336), .Y(n460) );
  CLKMX2X2 U448 ( .A(A[12]), .B(A[13]), .S0(n339), .Y(n470) );
  CLKMX2X2 U449 ( .A(A[14]), .B(A[15]), .S0(n339), .Y(n469) );
  MXI2X1 U450 ( .A(n471), .B(n403), .S0(n337), .Y(n387) );
  CLKMX2X2 U451 ( .A(A[8]), .B(A[9]), .S0(n339), .Y(n403) );
  CLKMX2X2 U452 ( .A(A[10]), .B(A[11]), .S0(n339), .Y(n471) );
endmodule


module alu_DW_leftsh_0 ( A, SH, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  wire   n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487;

  NAND4X1 U255 ( .A(n479), .B(n480), .C(n481), .D(n482), .Y(n321) );
  MXI3X1 U256 ( .A(n370), .B(n382), .C(n344), .S0(n339), .S1(n335), .Y(n322)
         );
  MXI3X1 U257 ( .A(n377), .B(n387), .C(n345), .S0(n339), .S1(n335), .Y(n323)
         );
  CLKINVX1 U258 ( .A(n391), .Y(n352) );
  CLKINVX1 U259 ( .A(n399), .Y(n347) );
  CLKINVX1 U260 ( .A(n393), .Y(n346) );
  INVX3 U261 ( .A(n340), .Y(n339) );
  INVX3 U262 ( .A(n336), .Y(n334) );
  INVX3 U263 ( .A(n340), .Y(n338) );
  INVX3 U264 ( .A(n336), .Y(n335) );
  INVX3 U265 ( .A(n333), .Y(n330) );
  INVX3 U266 ( .A(n332), .Y(n331) );
  CLKINVX1 U267 ( .A(n383), .Y(n344) );
  CLKINVX1 U268 ( .A(n388), .Y(n345) );
  CLKBUFX3 U269 ( .A(n337), .Y(n336) );
  CLKBUFX3 U270 ( .A(n341), .Y(n340) );
  CLKBUFX3 U271 ( .A(n325), .Y(n324) );
  INVX3 U272 ( .A(SH[0]), .Y(n343) );
  INVX3 U273 ( .A(SH[0]), .Y(n342) );
  CLKBUFX3 U274 ( .A(n333), .Y(n332) );
  CLKBUFX3 U275 ( .A(SH[4]), .Y(n329) );
  CLKBUFX3 U276 ( .A(SH[4]), .Y(n328) );
  CLKBUFX3 U277 ( .A(SH[5]), .Y(n327) );
  CLKBUFX3 U278 ( .A(SH[5]), .Y(n326) );
  CLKINVX1 U279 ( .A(n417), .Y(n348) );
  CLKINVX1 U280 ( .A(n422), .Y(n349) );
  CLKINVX1 U281 ( .A(n427), .Y(n350) );
  CLKINVX1 U282 ( .A(n432), .Y(n351) );
  CLKINVX1 U283 ( .A(n443), .Y(n353) );
  CLKINVX1 U284 ( .A(n403), .Y(n354) );
  CLKINVX1 U285 ( .A(n410), .Y(n355) );
  CLKINVX1 U286 ( .A(n363), .Y(n356) );
  CLKBUFX3 U287 ( .A(n321), .Y(n325) );
  CLKINVX1 U288 ( .A(SH[1]), .Y(n341) );
  CLKINVX1 U289 ( .A(SH[2]), .Y(n337) );
  CLKINVX1 U290 ( .A(SH[3]), .Y(n333) );
  NOR4X1 U291 ( .A(n326), .B(n329), .C(n357), .D(n325), .Y(B[9]) );
  NOR4X1 U292 ( .A(n326), .B(n328), .C(n358), .D(n321), .Y(B[8]) );
  NOR4X1 U293 ( .A(n327), .B(n328), .C(n325), .D(n359), .Y(B[7]) );
  NOR4X1 U294 ( .A(n327), .B(n328), .C(n325), .D(n360), .Y(B[6]) );
  NOR4X1 U295 ( .A(n327), .B(n328), .C(n325), .D(n361), .Y(B[5]) );
  NOR4X1 U296 ( .A(n326), .B(n328), .C(n325), .D(n362), .Y(B[4]) );
  NOR4X1 U297 ( .A(n327), .B(n329), .C(n321), .D(n363), .Y(B[3]) );
  NOR3X1 U298 ( .A(n364), .B(n327), .C(n325), .Y(B[31]) );
  MX3XL U299 ( .A(n365), .B(n366), .C(n367), .S0(n331), .S1(n328), .Y(n364) );
  MXI2X1 U300 ( .A(n368), .B(n369), .S0(n334), .Y(n365) );
  MX3XL U301 ( .A(A[31]), .B(A[30]), .C(n370), .S0(SH[0]), .S1(n339), .Y(n368)
         );
  NOR3X1 U302 ( .A(n371), .B(n327), .C(n325), .Y(B[30]) );
  MX3XL U303 ( .A(n372), .B(n373), .C(n374), .S0(n330), .S1(n328), .Y(n371) );
  MXI2X1 U304 ( .A(n375), .B(n376), .S0(n334), .Y(n372) );
  MX3XL U305 ( .A(A[30]), .B(A[29]), .C(n377), .S0(SH[0]), .S1(n339), .Y(n375)
         );
  NOR4X1 U306 ( .A(n326), .B(n329), .C(n325), .D(n378), .Y(B[2]) );
  NOR3X1 U307 ( .A(n379), .B(n327), .C(n324), .Y(B[29]) );
  MX3XL U308 ( .A(n322), .B(n380), .C(n381), .S0(n331), .S1(n328), .Y(n379) );
  CLKMX2X2 U309 ( .A(A[28]), .B(A[29]), .S0(n342), .Y(n370) );
  NOR3X1 U310 ( .A(n384), .B(n327), .C(n324), .Y(B[28]) );
  MX3XL U311 ( .A(n323), .B(n385), .C(n386), .S0(n331), .S1(n328), .Y(n384) );
  CLKMX2X2 U312 ( .A(A[27]), .B(A[28]), .S0(n342), .Y(n377) );
  NOR3X1 U313 ( .A(n389), .B(n327), .C(n324), .Y(B[27]) );
  MXI2X1 U314 ( .A(n390), .B(n352), .S0(n328), .Y(n389) );
  MX3XL U315 ( .A(n369), .B(n346), .C(n392), .S0(n335), .S1(n330), .Y(n390) );
  CLKMX2X2 U316 ( .A(n394), .B(n382), .S0(n340), .Y(n369) );
  CLKMX2X2 U317 ( .A(A[26]), .B(A[27]), .S0(n342), .Y(n382) );
  NOR3X1 U318 ( .A(n395), .B(n327), .C(n324), .Y(B[26]) );
  MX3XL U319 ( .A(n396), .B(n397), .C(n398), .S0(n331), .S1(n328), .Y(n395) );
  MXI2X1 U320 ( .A(n376), .B(n347), .S0(n335), .Y(n396) );
  CLKMX2X2 U321 ( .A(n400), .B(n387), .S0(n340), .Y(n376) );
  CLKMX2X2 U322 ( .A(A[25]), .B(A[26]), .S0(n342), .Y(n387) );
  NOR3X1 U323 ( .A(n401), .B(n327), .C(n324), .Y(B[25]) );
  CLKMX2X2 U324 ( .A(n402), .B(n357), .S0(n328), .Y(n401) );
  MXI2X1 U325 ( .A(n403), .B(n404), .S0(n330), .Y(n357) );
  MX3XL U326 ( .A(n383), .B(n405), .C(n406), .S0(n335), .S1(n330), .Y(n402) );
  MXI2X1 U327 ( .A(n394), .B(n407), .S0(n339), .Y(n383) );
  CLKMX2X2 U328 ( .A(A[24]), .B(A[25]), .S0(n342), .Y(n394) );
  NOR3X1 U329 ( .A(n408), .B(n327), .C(n324), .Y(B[24]) );
  CLKMX2X2 U330 ( .A(n409), .B(n358), .S0(n328), .Y(n408) );
  MXI2X1 U331 ( .A(n410), .B(n411), .S0(n330), .Y(n358) );
  MX3XL U332 ( .A(n388), .B(n412), .C(n413), .S0(n335), .S1(n330), .Y(n409) );
  MXI2X1 U333 ( .A(n400), .B(n414), .S0(n339), .Y(n388) );
  CLKMX2X2 U334 ( .A(A[23]), .B(A[24]), .S0(n342), .Y(n400) );
  NOR3X1 U335 ( .A(n415), .B(n327), .C(n324), .Y(B[23]) );
  MX3XL U336 ( .A(n366), .B(n348), .C(n359), .S0(n331), .S1(n328), .Y(n415) );
  NAND2X1 U337 ( .A(n416), .B(n332), .Y(n359) );
  CLKMX2X2 U338 ( .A(n418), .B(n393), .S0(n336), .Y(n366) );
  MXI2X1 U339 ( .A(n407), .B(n419), .S0(n339), .Y(n393) );
  CLKMX2X2 U340 ( .A(A[22]), .B(A[23]), .S0(n342), .Y(n407) );
  NOR3X1 U341 ( .A(n420), .B(n327), .C(n324), .Y(B[22]) );
  MX3XL U342 ( .A(n373), .B(n349), .C(n360), .S0(n331), .S1(n328), .Y(n420) );
  NAND2X1 U343 ( .A(n421), .B(n333), .Y(n360) );
  CLKMX2X2 U344 ( .A(n423), .B(n399), .S0(n336), .Y(n373) );
  MXI2X1 U345 ( .A(n414), .B(n424), .S0(n339), .Y(n399) );
  CLKMX2X2 U346 ( .A(A[21]), .B(A[22]), .S0(n342), .Y(n414) );
  NOR3X1 U347 ( .A(n425), .B(n327), .C(n324), .Y(B[21]) );
  MX3XL U348 ( .A(n380), .B(n350), .C(n361), .S0(n331), .S1(n328), .Y(n425) );
  NAND2X1 U349 ( .A(n426), .B(n333), .Y(n361) );
  CLKMX2X2 U350 ( .A(n428), .B(n405), .S0(n337), .Y(n380) );
  MXI2X1 U351 ( .A(n419), .B(n429), .S0(n339), .Y(n405) );
  CLKMX2X2 U352 ( .A(A[20]), .B(A[21]), .S0(n342), .Y(n419) );
  NOR3X1 U353 ( .A(n430), .B(n327), .C(n324), .Y(B[20]) );
  MX3XL U354 ( .A(n385), .B(n351), .C(n362), .S0(n331), .S1(n329), .Y(n430) );
  NAND2X1 U355 ( .A(n431), .B(n333), .Y(n362) );
  CLKMX2X2 U356 ( .A(n433), .B(n412), .S0(n336), .Y(n385) );
  MXI2X1 U357 ( .A(n424), .B(n434), .S0(n339), .Y(n412) );
  CLKMX2X2 U358 ( .A(A[19]), .B(A[20]), .S0(n342), .Y(n424) );
  NOR4X1 U359 ( .A(n326), .B(n329), .C(n321), .D(n435), .Y(B[1]) );
  NOR3BXL U360 ( .AN(n436), .B(n327), .C(n325), .Y(B[19]) );
  MX3XL U361 ( .A(n392), .B(n437), .C(n356), .S0(n331), .S1(n329), .Y(n436) );
  NAND2X1 U362 ( .A(n438), .B(n332), .Y(n363) );
  MXI2X1 U363 ( .A(n418), .B(n439), .S0(n335), .Y(n392) );
  MXI2X1 U364 ( .A(n429), .B(n440), .S0(n339), .Y(n418) );
  CLKMX2X2 U365 ( .A(A[18]), .B(A[19]), .S0(n342), .Y(n429) );
  NOR3X1 U366 ( .A(n441), .B(SH[5]), .C(n325), .Y(B[18]) );
  MX3XL U367 ( .A(n397), .B(n353), .C(n378), .S0(n331), .S1(n328), .Y(n441) );
  NAND2X1 U368 ( .A(n442), .B(n333), .Y(n378) );
  CLKMX2X2 U369 ( .A(n444), .B(n423), .S0(n336), .Y(n397) );
  MXI2X1 U370 ( .A(n434), .B(n445), .S0(n339), .Y(n423) );
  CLKMX2X2 U371 ( .A(A[17]), .B(A[18]), .S0(n342), .Y(n434) );
  NOR3X1 U372 ( .A(n446), .B(SH[5]), .C(n325), .Y(B[17]) );
  MX3XL U373 ( .A(n406), .B(n354), .C(n435), .S0(n331), .S1(n329), .Y(n446) );
  NAND2X1 U374 ( .A(n404), .B(n332), .Y(n435) );
  NOR2X1 U375 ( .A(n447), .B(n335), .Y(n404) );
  MXI2X1 U376 ( .A(n448), .B(n449), .S0(n335), .Y(n403) );
  CLKMX2X2 U377 ( .A(n450), .B(n428), .S0(n336), .Y(n406) );
  MXI2X1 U378 ( .A(n440), .B(n451), .S0(n339), .Y(n428) );
  CLKMX2X2 U379 ( .A(A[16]), .B(A[17]), .S0(n342), .Y(n440) );
  NOR3X1 U380 ( .A(n452), .B(SH[5]), .C(n325), .Y(B[16]) );
  MX3XL U381 ( .A(n413), .B(n355), .C(n453), .S0(n330), .S1(n328), .Y(n452) );
  MXI2X1 U382 ( .A(n454), .B(n455), .S0(n334), .Y(n410) );
  CLKMX2X2 U383 ( .A(n456), .B(n433), .S0(n336), .Y(n413) );
  MXI2X1 U384 ( .A(n445), .B(n457), .S0(n339), .Y(n433) );
  CLKMX2X2 U385 ( .A(A[15]), .B(A[16]), .S0(n343), .Y(n445) );
  NOR4X1 U386 ( .A(n326), .B(n329), .C(n367), .D(n325), .Y(B[15]) );
  MXI2X1 U387 ( .A(n417), .B(n416), .S0(n330), .Y(n367) );
  MXI2X1 U388 ( .A(n458), .B(n459), .S0(n334), .Y(n416) );
  MXI2X1 U389 ( .A(n439), .B(n460), .S0(n334), .Y(n417) );
  MXI2X1 U390 ( .A(n451), .B(n461), .S0(n338), .Y(n439) );
  CLKMX2X2 U391 ( .A(A[14]), .B(A[15]), .S0(n343), .Y(n451) );
  NOR4X1 U392 ( .A(n326), .B(n329), .C(n374), .D(n324), .Y(B[14]) );
  MXI2X1 U393 ( .A(n422), .B(n421), .S0(n330), .Y(n374) );
  MXI2X1 U394 ( .A(n462), .B(n463), .S0(n334), .Y(n421) );
  MXI2X1 U395 ( .A(n444), .B(n464), .S0(n334), .Y(n422) );
  MXI2X1 U396 ( .A(n457), .B(n465), .S0(n338), .Y(n444) );
  CLKMX2X2 U397 ( .A(A[13]), .B(A[14]), .S0(n343), .Y(n457) );
  NOR4X1 U398 ( .A(n326), .B(n329), .C(n381), .D(n324), .Y(B[13]) );
  MXI2X1 U399 ( .A(n427), .B(n426), .S0(n330), .Y(n381) );
  MXI2X1 U400 ( .A(n449), .B(n447), .S0(n334), .Y(n426) );
  NAND2X1 U401 ( .A(n466), .B(n340), .Y(n447) );
  MXI2X1 U402 ( .A(n467), .B(n468), .S0(n338), .Y(n449) );
  MXI2X1 U403 ( .A(n450), .B(n448), .S0(n334), .Y(n427) );
  MXI2X1 U404 ( .A(n469), .B(n470), .S0(n338), .Y(n448) );
  MXI2X1 U405 ( .A(n461), .B(n471), .S0(n338), .Y(n450) );
  CLKMX2X2 U406 ( .A(A[12]), .B(A[13]), .S0(n343), .Y(n461) );
  NOR4X1 U407 ( .A(n326), .B(n329), .C(n386), .D(n324), .Y(B[12]) );
  MXI2X1 U408 ( .A(n432), .B(n431), .S0(n330), .Y(n386) );
  MXI2X1 U409 ( .A(n455), .B(n472), .S0(n334), .Y(n431) );
  MXI2X1 U410 ( .A(n473), .B(n474), .S0(n338), .Y(n455) );
  MXI2X1 U411 ( .A(n456), .B(n454), .S0(n334), .Y(n432) );
  MXI2X1 U412 ( .A(n475), .B(n476), .S0(n338), .Y(n454) );
  MXI2X1 U413 ( .A(n465), .B(n477), .S0(n338), .Y(n456) );
  CLKMX2X2 U414 ( .A(A[11]), .B(A[12]), .S0(n343), .Y(n465) );
  NOR4X1 U415 ( .A(n326), .B(n329), .C(n391), .D(n321), .Y(B[11]) );
  MXI2X1 U416 ( .A(n437), .B(n438), .S0(n330), .Y(n391) );
  NOR2X1 U417 ( .A(n459), .B(n335), .Y(n438) );
  MXI2X1 U418 ( .A(n468), .B(n466), .S0(n338), .Y(n459) );
  CLKMX2X2 U419 ( .A(A[0]), .B(A[1]), .S0(n343), .Y(n466) );
  CLKMX2X2 U420 ( .A(A[2]), .B(A[3]), .S0(n343), .Y(n468) );
  MXI2X1 U421 ( .A(n460), .B(n458), .S0(n334), .Y(n437) );
  MXI2X1 U422 ( .A(n470), .B(n467), .S0(n338), .Y(n458) );
  CLKMX2X2 U423 ( .A(A[4]), .B(A[5]), .S0(n343), .Y(n467) );
  CLKMX2X2 U424 ( .A(A[6]), .B(A[7]), .S0(n343), .Y(n470) );
  MXI2X1 U425 ( .A(n471), .B(n469), .S0(n338), .Y(n460) );
  CLKMX2X2 U426 ( .A(A[8]), .B(A[9]), .S0(n343), .Y(n469) );
  CLKMX2X2 U427 ( .A(A[10]), .B(A[11]), .S0(n343), .Y(n471) );
  NOR4X1 U428 ( .A(n326), .B(n329), .C(n398), .D(n325), .Y(B[10]) );
  MXI2X1 U429 ( .A(n443), .B(n442), .S0(n330), .Y(n398) );
  NOR2X1 U430 ( .A(n463), .B(n335), .Y(n442) );
  MXI2X1 U431 ( .A(n474), .B(n478), .S0(n338), .Y(n463) );
  CLKMX2X2 U432 ( .A(A[1]), .B(A[2]), .S0(n343), .Y(n474) );
  MXI2X1 U433 ( .A(n464), .B(n462), .S0(n334), .Y(n443) );
  MXI2X1 U434 ( .A(n476), .B(n473), .S0(n338), .Y(n462) );
  CLKMX2X2 U435 ( .A(A[3]), .B(A[4]), .S0(n343), .Y(n473) );
  CLKMX2X2 U436 ( .A(A[5]), .B(A[6]), .S0(n342), .Y(n476) );
  MXI2X1 U437 ( .A(n477), .B(n475), .S0(n339), .Y(n464) );
  CLKMX2X2 U438 ( .A(A[7]), .B(A[8]), .S0(n342), .Y(n475) );
  CLKMX2X2 U439 ( .A(A[9]), .B(A[10]), .S0(n342), .Y(n477) );
  NOR4X1 U440 ( .A(n326), .B(n329), .C(n321), .D(n453), .Y(B[0]) );
  NAND2X1 U441 ( .A(n411), .B(n332), .Y(n453) );
  NOR2X1 U442 ( .A(n472), .B(n335), .Y(n411) );
  NAND2X1 U443 ( .A(n478), .B(n340), .Y(n472) );
  NOR2BX1 U444 ( .AN(A[0]), .B(SH[0]), .Y(n478) );
  AND4X1 U445 ( .A(n483), .B(n484), .C(n485), .D(n486), .Y(n482) );
  NOR4X1 U446 ( .A(SH[9]), .B(SH[8]), .C(SH[7]), .D(SH[6]), .Y(n486) );
  NOR3X1 U447 ( .A(SH[29]), .B(SH[31]), .C(SH[30]), .Y(n485) );
  NOR3X1 U448 ( .A(SH[26]), .B(SH[28]), .C(SH[27]), .Y(n484) );
  NOR3X1 U449 ( .A(SH[23]), .B(SH[25]), .C(SH[24]), .Y(n483) );
  NOR4X1 U450 ( .A(n487), .B(SH[16]), .C(SH[18]), .D(SH[17]), .Y(n481) );
  OR4X1 U451 ( .A(SH[20]), .B(SH[19]), .C(SH[22]), .D(SH[21]), .Y(n487) );
  NOR3X1 U452 ( .A(SH[13]), .B(SH[15]), .C(SH[14]), .Y(n480) );
  NOR3X1 U453 ( .A(SH[10]), .B(SH[12]), .C(SH[11]), .Y(n479) );
endmodule


module alu_DW_cmp_0 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375;

  CLKINVX1 U655 ( .A(A[1]), .Y(n1281) );
  OAI2BB1X1 U656 ( .A0N(n1332), .A1N(n1278), .B0(n1321), .Y(n1319) );
  OA22X1 U657 ( .A0(n1327), .A1(n1328), .B0(n1329), .B1(n1327), .Y(n1278) );
  CLKINVX1 U658 ( .A(B[3]), .Y(n1312) );
  CLKINVX1 U659 ( .A(B[2]), .Y(n1313) );
  CLKINVX1 U660 ( .A(B[24]), .Y(n1290) );
  CLKINVX1 U661 ( .A(B[18]), .Y(n1297) );
  CLKINVX1 U662 ( .A(B[14]), .Y(n1301) );
  CLKINVX1 U663 ( .A(B[26]), .Y(n1288) );
  CLKINVX1 U664 ( .A(B[20]), .Y(n1295) );
  CLKINVX1 U665 ( .A(B[22]), .Y(n1293) );
  CLKINVX1 U666 ( .A(B[30]), .Y(n1283) );
  CLKINVX1 U667 ( .A(B[16]), .Y(n1299) );
  CLKINVX1 U668 ( .A(B[6]), .Y(n1311) );
  CLKINVX1 U669 ( .A(B[17]), .Y(n1298) );
  CLKINVX1 U670 ( .A(B[15]), .Y(n1300) );
  CLKINVX1 U671 ( .A(B[7]), .Y(n1310) );
  CLKINVX1 U672 ( .A(B[31]), .Y(n1282) );
  CLKINVX1 U673 ( .A(n1338), .Y(n1284) );
  CLKINVX1 U674 ( .A(A[4]), .Y(n1280) );
  CLKINVX1 U675 ( .A(A[5]), .Y(n1279) );
  CLKINVX1 U676 ( .A(n1324), .Y(n1292) );
  CLKINVX1 U677 ( .A(B[19]), .Y(n1296) );
  CLKINVX1 U678 ( .A(B[23]), .Y(n1291) );
  CLKINVX1 U679 ( .A(B[27]), .Y(n1287) );
  CLKINVX1 U680 ( .A(n1369), .Y(n1302) );
  CLKINVX1 U681 ( .A(B[21]), .Y(n1294) );
  CLKINVX1 U682 ( .A(B[25]), .Y(n1289) );
  CLKINVX1 U683 ( .A(n1359), .Y(n1309) );
  CLKINVX1 U684 ( .A(A[12]), .Y(n1304) );
  CLKINVX1 U685 ( .A(A[28]), .Y(n1286) );
  CLKINVX1 U686 ( .A(A[8]), .Y(n1308) );
  CLKINVX1 U687 ( .A(A[10]), .Y(n1306) );
  CLKINVX1 U688 ( .A(A[9]), .Y(n1307) );
  CLKINVX1 U689 ( .A(A[11]), .Y(n1305) );
  CLKINVX1 U690 ( .A(A[29]), .Y(n1285) );
  CLKINVX1 U691 ( .A(A[13]), .Y(n1303) );
  OAI31XL U692 ( .A0(n1314), .A1(n1315), .A2(n1316), .B0(n1317), .Y(
        GE_LT_GT_LE) );
  OAI22XL U693 ( .A0(n1318), .A1(n1319), .B0(n1320), .B1(n1318), .Y(n1317) );
  OAI22XL U694 ( .A0(n1322), .A1(n1323), .B0(n1324), .B1(n1322), .Y(n1321) );
  OAI32X1 U695 ( .A0(n1295), .A1(A[20]), .A2(n1325), .B0(A[21]), .B1(n1294), 
        .Y(n1323) );
  OAI32X1 U696 ( .A0(n1293), .A1(A[22]), .A2(n1326), .B0(A[23]), .B1(n1291), 
        .Y(n1322) );
  OAI32X1 U697 ( .A0(n1299), .A1(A[16]), .A2(n1330), .B0(A[17]), .B1(n1298), 
        .Y(n1328) );
  OAI32X1 U698 ( .A0(n1297), .A1(A[18]), .A2(n1331), .B0(A[19]), .B1(n1296), 
        .Y(n1327) );
  OAI21XL U699 ( .A0(n1333), .A1(n1334), .B0(n1335), .Y(n1318) );
  OAI22XL U700 ( .A0(n1336), .A1(n1284), .B0(n1337), .B1(n1336), .Y(n1335) );
  AOI32X1 U701 ( .A0(B[28]), .A1(n1286), .A2(n1339), .B0(n1285), .B1(B[29]), 
        .Y(n1338) );
  OAI32X1 U702 ( .A0(n1283), .A1(A[30]), .A2(n1340), .B0(A[31]), .B1(n1282), 
        .Y(n1336) );
  OAI22XL U703 ( .A0(n1341), .A1(n1342), .B0(n1343), .B1(n1341), .Y(n1334) );
  OAI32X1 U704 ( .A0(n1290), .A1(A[24]), .A2(n1344), .B0(A[25]), .B1(n1289), 
        .Y(n1342) );
  OAI32X1 U705 ( .A0(n1288), .A1(A[26]), .A2(n1345), .B0(A[27]), .B1(n1287), 
        .Y(n1341) );
  OAI22XL U706 ( .A0(n1346), .A1(n1347), .B0(n1348), .B1(n1346), .Y(n1316) );
  NOR3X1 U707 ( .A(n1349), .B(n1350), .C(n1351), .Y(n1348) );
  OAI21XL U708 ( .A0(B[8]), .A1(n1308), .B0(n1352), .Y(n1349) );
  OAI31XL U709 ( .A0(n1353), .A1(n1354), .A2(n1355), .B0(n1356), .Y(n1347) );
  AO22X1 U710 ( .A0(n1309), .A1(n1357), .B0(n1355), .B1(n1309), .Y(n1356) );
  AOI32X1 U711 ( .A0(B[4]), .A1(n1280), .A2(n1358), .B0(n1279), .B1(B[5]), .Y(
        n1357) );
  OAI32X1 U712 ( .A0(n1311), .A1(A[6]), .A2(n1360), .B0(A[7]), .B1(n1310), .Y(
        n1359) );
  AO21X1 U713 ( .A0(n1311), .A1(A[6]), .B0(n1360), .Y(n1355) );
  NOR2BX1 U714 ( .AN(A[7]), .B(B[7]), .Y(n1360) );
  AOI221XL U715 ( .A0(B[1]), .A1(n1281), .B0(n1361), .B1(B[0]), .C0(n1362), 
        .Y(n1354) );
  AOI2BB1X1 U716 ( .A0N(n1281), .A1N(B[1]), .B0(A[0]), .Y(n1361) );
  OAI221XL U717 ( .A0(B[4]), .A1(n1280), .B0(n1363), .B1(n1362), .C0(n1358), 
        .Y(n1353) );
  OR2X1 U718 ( .A(B[5]), .B(n1279), .Y(n1358) );
  OAI32X1 U719 ( .A0(n1313), .A1(A[2]), .A2(n1364), .B0(A[3]), .B1(n1312), .Y(
        n1362) );
  AOI21X1 U720 ( .A0(A[2]), .A1(n1313), .B0(n1364), .Y(n1363) );
  AND2X1 U721 ( .A(A[3]), .B(n1312), .Y(n1364) );
  OAI21XL U722 ( .A0(n1350), .A1(n1365), .B0(n1366), .Y(n1346) );
  OAI22XL U723 ( .A0(n1367), .A1(n1302), .B0(n1368), .B1(n1367), .Y(n1366) );
  AOI32X1 U724 ( .A0(B[12]), .A1(n1304), .A2(n1370), .B0(n1303), .B1(B[13]), 
        .Y(n1369) );
  OAI32X1 U725 ( .A0(n1301), .A1(A[14]), .A2(n1371), .B0(A[15]), .B1(n1300), 
        .Y(n1367) );
  AO22X1 U726 ( .A0(n1372), .A1(n1373), .B0(n1351), .B1(n1372), .Y(n1365) );
  OAI21XL U727 ( .A0(B[10]), .A1(n1306), .B0(n1374), .Y(n1351) );
  AOI32X1 U728 ( .A0(B[8]), .A1(n1308), .A2(n1352), .B0(n1307), .B1(B[9]), .Y(
        n1373) );
  OR2X1 U729 ( .A(B[9]), .B(n1307), .Y(n1352) );
  AOI32X1 U730 ( .A0(B[10]), .A1(n1306), .A2(n1374), .B0(n1305), .B1(B[11]), 
        .Y(n1372) );
  OR2X1 U731 ( .A(B[11]), .B(n1305), .Y(n1374) );
  OAI211X1 U732 ( .A0(B[12]), .A1(n1304), .B0(n1370), .C0(n1368), .Y(n1350) );
  AOI21X1 U733 ( .A0(n1301), .A1(A[14]), .B0(n1371), .Y(n1368) );
  NOR2BX1 U734 ( .AN(A[15]), .B(B[15]), .Y(n1371) );
  OR2X1 U735 ( .A(B[13]), .B(n1303), .Y(n1370) );
  AO21X1 U736 ( .A0(n1299), .A1(A[16]), .B0(n1330), .Y(n1315) );
  AND2X1 U737 ( .A(A[17]), .B(n1298), .Y(n1330) );
  NAND3X1 U738 ( .A(n1320), .B(n1332), .C(n1329), .Y(n1314) );
  AOI21X1 U739 ( .A0(n1297), .A1(A[18]), .B0(n1331), .Y(n1329) );
  NOR2BX1 U740 ( .AN(A[19]), .B(B[19]), .Y(n1331) );
  AOI211X1 U741 ( .A0(n1295), .A1(A[20]), .B0(n1325), .C0(n1292), .Y(n1332) );
  AOI21X1 U742 ( .A0(n1293), .A1(A[22]), .B0(n1326), .Y(n1324) );
  NOR2BX1 U743 ( .AN(A[23]), .B(B[23]), .Y(n1326) );
  NOR2BX1 U744 ( .AN(A[21]), .B(B[21]), .Y(n1325) );
  AOI211X1 U745 ( .A0(n1290), .A1(A[24]), .B0(n1344), .C0(n1375), .Y(n1320) );
  NAND2BX1 U746 ( .AN(n1333), .B(n1343), .Y(n1375) );
  AOI21X1 U747 ( .A0(n1288), .A1(A[26]), .B0(n1345), .Y(n1343) );
  NOR2BX1 U748 ( .AN(A[27]), .B(B[27]), .Y(n1345) );
  OAI211X1 U749 ( .A0(B[28]), .A1(n1286), .B0(n1339), .C0(n1337), .Y(n1333) );
  AOI21X1 U750 ( .A0(n1283), .A1(A[30]), .B0(n1340), .Y(n1337) );
  NOR2BX1 U751 ( .AN(A[31]), .B(B[31]), .Y(n1340) );
  OR2X1 U752 ( .A(B[29]), .B(n1285), .Y(n1339) );
  NOR2BX1 U753 ( .AN(A[25]), .B(B[25]), .Y(n1344) );
endmodule


module alu_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [32:0] carry;

  ADDFXL U2_30 ( .A(A[30]), .B(n6), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  ADDFXL U2_29 ( .A(A[29]), .B(n7), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  ADDFXL U2_26 ( .A(A[26]), .B(n10), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  ADDFXL U2_24 ( .A(A[24]), .B(n12), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  ADDFXL U2_22 ( .A(A[22]), .B(n14), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  ADDFXL U2_20 ( .A(A[20]), .B(n16), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  ADDFXL U2_18 ( .A(A[18]), .B(n18), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  ADDFXL U2_17 ( .A(A[17]), .B(n19), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  ADDFXL U2_16 ( .A(A[16]), .B(n20), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n22), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_6 ( .A(A[6]), .B(n30), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_28 ( .A(A[28]), .B(n8), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n23), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n24), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n25), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n26), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n27), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n28), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  ADDFXL U2_27 ( .A(A[27]), .B(n9), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  ADDFXL U2_25 ( .A(A[25]), .B(n11), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  ADDFXL U2_23 ( .A(A[23]), .B(n13), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  ADDFXL U2_21 ( .A(A[21]), .B(n15), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  ADDFXL U2_19 ( .A(A[19]), .B(n17), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  ADDFXL U2_15 ( .A(A[15]), .B(n21), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  ADDFXL U2_7 ( .A(A[7]), .B(n29), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  XOR3X1 U2_31 ( .A(A[31]), .B(n5), .C(carry[31]), .Y(DIFF[31]) );
  ADDFXL U2_5 ( .A(A[5]), .B(n4), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADDFXL U2_4 ( .A(A[4]), .B(n3), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADDFXL U2_2 ( .A(A[2]), .B(n32), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n33), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n31), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  CLKINVX1 U1 ( .A(B[0]), .Y(n2) );
  CLKINVX1 U2 ( .A(B[3]), .Y(n31) );
  NAND2X1 U3 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U4 ( .A(B[1]), .Y(n33) );
  CLKINVX1 U5 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U6 ( .A(B[2]), .Y(n32) );
  CLKINVX1 U7 ( .A(B[4]), .Y(n3) );
  CLKINVX1 U8 ( .A(B[5]), .Y(n4) );
  XNOR2X1 U9 ( .A(n2), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U10 ( .A(B[31]), .Y(n5) );
  CLKINVX1 U11 ( .A(B[7]), .Y(n29) );
  CLKINVX1 U12 ( .A(B[15]), .Y(n21) );
  CLKINVX1 U13 ( .A(B[19]), .Y(n17) );
  CLKINVX1 U14 ( .A(B[21]), .Y(n15) );
  CLKINVX1 U15 ( .A(B[23]), .Y(n13) );
  CLKINVX1 U16 ( .A(B[25]), .Y(n11) );
  CLKINVX1 U17 ( .A(B[27]), .Y(n9) );
  CLKINVX1 U18 ( .A(B[8]), .Y(n28) );
  CLKINVX1 U19 ( .A(B[9]), .Y(n27) );
  CLKINVX1 U20 ( .A(B[10]), .Y(n26) );
  CLKINVX1 U21 ( .A(B[11]), .Y(n25) );
  CLKINVX1 U22 ( .A(B[12]), .Y(n24) );
  CLKINVX1 U23 ( .A(B[13]), .Y(n23) );
  CLKINVX1 U24 ( .A(B[28]), .Y(n8) );
  CLKINVX1 U25 ( .A(B[6]), .Y(n30) );
  CLKINVX1 U26 ( .A(B[14]), .Y(n22) );
  CLKINVX1 U27 ( .A(B[16]), .Y(n20) );
  CLKINVX1 U28 ( .A(B[17]), .Y(n19) );
  CLKINVX1 U29 ( .A(B[18]), .Y(n18) );
  CLKINVX1 U30 ( .A(B[20]), .Y(n16) );
  CLKINVX1 U31 ( .A(B[22]), .Y(n14) );
  CLKINVX1 U32 ( .A(B[24]), .Y(n12) );
  CLKINVX1 U33 ( .A(B[26]), .Y(n10) );
  CLKINVX1 U34 ( .A(B[29]), .Y(n7) );
  CLKINVX1 U35 ( .A(B[30]), .Y(n6) );
endmodule


module alu_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  XOR3X1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module alu ( ctrl, x, y, out );
  input [3:0] ctrl;
  input [31:0] x;
  input [31:0] y;
  output [31:0] out;
  wire   N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72,
         N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N205, N206, N207,
         N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218,
         N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251,
         N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262,
         N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273,
         N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284,
         N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295,
         N296, N297, N298, N299, N300, N301, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301;

  alu_DW_rightsh_0 srl_179 ( .A({n32, n31, n30, n29, n28, n27, n26, n25, n24, 
        n23, n22, n21, n20, n19, n12, n11, n10, n9, n8, n7, n6, n5, n4, n3, n2, 
        n1, n53, n260, n262, n264, n266, n268}), .DATA_TC(1'b0), .SH({y[31:6], 
        n273, n272, y[3:1], n270}), .B({N301, N300, N299, N298, N297, N296, 
        N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, 
        N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, 
        N271, N270}) );
  alu_DW_rightsh_1 sra_176 ( .A({y[31:6], n273, n272, y[3:1], n270}), 
        .DATA_TC(1'b0), .SH({n32, n31, n30, n29, n28, n27, n26, n25, n24, n23, 
        n22, n21, n20, n19, n12, n11, n10, n9, n8, n7, n6, n5, n4, n3, n2, n1, 
        n53, n260, n262, n264, n266, n268}), .B({N269, N268, N267, N266, N265, 
        N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, 
        N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, 
        N240, N239, N238}) );
  alu_DW_leftsh_0 sll_173 ( .A({y[31:6], n273, n272, y[3:1], n270}), .SH({n32, 
        n31, n30, n29, n28, n27, n26, n25, n24, n23, n22, n21, n20, n19, n12, 
        n11, n10, n9, n8, n7, n6, n5, n4, n3, n2, n1, n53, n260, n262, n264, 
        n266, n268}), .B({N237, N236, N235, N234, N233, N232, N231, N230, N229, 
        N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, 
        N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206}) );
  alu_DW_cmp_0 lt_166 ( .A({n32, n31, n30, n29, n28, n27, n26, n25, n24, n23, 
        n22, n21, n20, n19, n12, n11, n10, n9, n8, n7, n6, n5, n4, n3, n2, n1, 
        n53, n260, n262, n264, n266, n268}), .B({y[31:6], n273, n272, y[3:1], 
        n270}), .TC(1'b0), .GE_LT(1'b1), .GE_GT_EQ(1'b0), .GE_LT_GT_LE(N205)
         );
  alu_DW01_sub_0 sub_151 ( .A({n32, n31, n30, n29, n28, n27, n26, n25, n24, 
        n23, n22, n21, n20, n19, n12, n11, n10, n9, n8, n7, n6, n5, n4, n3, n2, 
        n1, n53, n260, n262, n264, n266, n268}), .B({y[31:6], n273, n272, 
        y[3:1], n270}), .CI(1'b0), .DIFF({N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77}) );
  alu_DW01_add_0 add_148 ( .A({n32, n31, n30, n29, n28, n27, n26, n25, n24, 
        n23, n22, n21, n20, n19, n12, n11, n10, n9, n8, n7, n6, n5, n4, n3, n2, 
        n1, n53, n260, n262, n264, n266, n268}), .B({y[31:6], n273, n272, 
        y[3:1], n270}), .CI(1'b0), .SUM({N76, N75, N74, N73, N72, N71, N70, 
        N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45}) );
  CLKBUFX3 U5 ( .A(n67), .Y(n35) );
  NAND2X1 U6 ( .A(n254), .B(n300), .Y(n66) );
  INVX3 U7 ( .A(n269), .Y(n268) );
  INVX3 U8 ( .A(n267), .Y(n266) );
  CLKINVX1 U9 ( .A(y[0]), .Y(n271) );
  CLKBUFX3 U10 ( .A(y[5]), .Y(n273) );
  CLKBUFX3 U14 ( .A(y[4]), .Y(n272) );
  INVX3 U15 ( .A(n263), .Y(n262) );
  INVX3 U16 ( .A(n261), .Y(n260) );
  INVX3 U17 ( .A(n259), .Y(n53) );
  CLKINVX1 U18 ( .A(x[0]), .Y(n269) );
  CLKINVX1 U19 ( .A(x[2]), .Y(n265) );
  CLKINVX1 U20 ( .A(x[1]), .Y(n267) );
  CLKINVX1 U21 ( .A(x[4]), .Y(n261) );
  CLKINVX1 U22 ( .A(x[3]), .Y(n263) );
  CLKINVX1 U23 ( .A(x[5]), .Y(n259) );
  AOI22X1 U24 ( .A0(N293), .A1(n35), .B0(N261), .B1(n34), .Y(n161) );
  AOI22X1 U25 ( .A0(N292), .A1(n35), .B0(N260), .B1(n34), .Y(n167) );
  AOI22X1 U26 ( .A0(N279), .A1(n36), .B0(N247), .B1(n68), .Y(n54) );
  AOI22X1 U27 ( .A0(N291), .A1(n35), .B0(N259), .B1(n34), .Y(n173) );
  AOI22X1 U28 ( .A0(N285), .A1(n36), .B0(N253), .B1(n33), .Y(n215) );
  AOI22X1 U29 ( .A0(N284), .A1(n67), .B0(N252), .B1(n33), .Y(n221) );
  AOI22X1 U30 ( .A0(N283), .A1(n67), .B0(N251), .B1(n33), .Y(n227) );
  AOI22X1 U31 ( .A0(N281), .A1(n67), .B0(N249), .B1(n33), .Y(n239) );
  AOI22X1 U32 ( .A0(N280), .A1(n67), .B0(N248), .B1(n33), .Y(n245) );
  AOI22X1 U33 ( .A0(N272), .A1(n35), .B0(N240), .B1(n34), .Y(n119) );
  CLKBUFX3 U34 ( .A(n60), .Y(n48) );
  CLKBUFX3 U35 ( .A(n68), .Y(n33) );
  CLKBUFX3 U36 ( .A(n68), .Y(n34) );
  CLKBUFX3 U37 ( .A(n60), .Y(n47) );
  CLKBUFX3 U38 ( .A(n60), .Y(n46) );
  CLKBUFX3 U39 ( .A(n64), .Y(n43) );
  CLKBUFX3 U40 ( .A(n64), .Y(n41) );
  CLKBUFX3 U41 ( .A(n65), .Y(n39) );
  CLKBUFX3 U42 ( .A(n64), .Y(n42) );
  CLKBUFX3 U43 ( .A(n66), .Y(n37) );
  CLKBUFX3 U44 ( .A(n66), .Y(n38) );
  CLKBUFX3 U45 ( .A(n65), .Y(n40) );
  AOI22X1 U46 ( .A0(N290), .A1(n35), .B0(N258), .B1(n33), .Y(n179) );
  AOI22X1 U47 ( .A0(N282), .A1(n67), .B0(N250), .B1(n33), .Y(n233) );
  AOI22X1 U48 ( .A0(N270), .A1(n67), .B0(N238), .B1(n33), .Y(n249) );
  AOI22X1 U49 ( .A0(N300), .A1(n35), .B0(N268), .B1(n34), .Y(n113) );
  AOI22X1 U50 ( .A0(N299), .A1(n35), .B0(N267), .B1(n34), .Y(n125) );
  AOI22X1 U51 ( .A0(N298), .A1(n35), .B0(N266), .B1(n34), .Y(n131) );
  AOI22X1 U52 ( .A0(N297), .A1(n35), .B0(N265), .B1(n34), .Y(n137) );
  AOI22X1 U53 ( .A0(N296), .A1(n35), .B0(N264), .B1(n34), .Y(n143) );
  AOI22X1 U54 ( .A0(N295), .A1(n35), .B0(N263), .B1(n34), .Y(n149) );
  AOI22X1 U55 ( .A0(N294), .A1(n35), .B0(N262), .B1(n34), .Y(n155) );
  AOI22X1 U56 ( .A0(N289), .A1(n36), .B0(N257), .B1(n33), .Y(n191) );
  AOI22X1 U57 ( .A0(N288), .A1(n36), .B0(N256), .B1(n33), .Y(n197) );
  AOI22X1 U58 ( .A0(N287), .A1(n36), .B0(N255), .B1(n33), .Y(n203) );
  AOI22X1 U59 ( .A0(N286), .A1(n36), .B0(N254), .B1(n33), .Y(n209) );
  AOI22X1 U60 ( .A0(N273), .A1(n36), .B0(N241), .B1(n34), .Y(n101) );
  AOI22X1 U61 ( .A0(N271), .A1(n35), .B0(N239), .B1(n33), .Y(n185) );
  AOI22X1 U62 ( .A0(N301), .A1(n36), .B0(N269), .B1(n34), .Y(n107) );
  AOI22X1 U63 ( .A0(N278), .A1(n36), .B0(N246), .B1(n34), .Y(n71) );
  AOI22X1 U64 ( .A0(N277), .A1(n36), .B0(N245), .B1(n33), .Y(n77) );
  AOI22X1 U65 ( .A0(N276), .A1(n36), .B0(N244), .B1(n68), .Y(n83) );
  AOI22X1 U66 ( .A0(N275), .A1(n36), .B0(N243), .B1(n68), .Y(n89) );
  AOI22X1 U67 ( .A0(N274), .A1(n36), .B0(N242), .B1(n68), .Y(n95) );
  AND2X2 U68 ( .A(n258), .B(n301), .Y(n68) );
  AOI22X1 U69 ( .A0(N82), .A1(n51), .B0(N50), .B1(n49), .Y(n87) );
  AOI22X1 U70 ( .A0(N81), .A1(n51), .B0(N49), .B1(n49), .Y(n93) );
  AOI22X1 U71 ( .A0(N80), .A1(n51), .B0(N48), .B1(n49), .Y(n99) );
  AOI22X1 U72 ( .A0(N79), .A1(n51), .B0(N47), .B1(n49), .Y(n117) );
  NAND3X1 U73 ( .A(n301), .B(n300), .C(n253), .Y(n65) );
  CLKBUFX3 U74 ( .A(n58), .Y(n50) );
  CLKBUFX3 U75 ( .A(n58), .Y(n49) );
  CLKBUFX3 U76 ( .A(n57), .Y(n51) );
  CLKBUFX3 U77 ( .A(n61), .Y(n45) );
  CLKBUFX3 U78 ( .A(n61), .Y(n44) );
  CLKBUFX3 U79 ( .A(n67), .Y(n36) );
  CLKBUFX3 U80 ( .A(n57), .Y(n52) );
  AOI22X1 U81 ( .A0(N107), .A1(n51), .B0(N75), .B1(n50), .Y(n111) );
  AOI22X1 U82 ( .A0(N106), .A1(n51), .B0(N74), .B1(n49), .Y(n123) );
  AOI22X1 U83 ( .A0(N105), .A1(n51), .B0(N73), .B1(n49), .Y(n129) );
  AOI22X1 U84 ( .A0(N104), .A1(n51), .B0(N72), .B1(n49), .Y(n135) );
  AOI22X1 U85 ( .A0(N103), .A1(n51), .B0(N71), .B1(n49), .Y(n141) );
  AOI22X1 U86 ( .A0(N102), .A1(n57), .B0(N70), .B1(n49), .Y(n147) );
  AOI22X1 U87 ( .A0(N101), .A1(n57), .B0(N69), .B1(n50), .Y(n153) );
  AOI22X1 U88 ( .A0(N100), .A1(n57), .B0(N68), .B1(n50), .Y(n159) );
  INVX3 U89 ( .A(n271), .Y(n270) );
  AOI22X1 U90 ( .A0(N99), .A1(n52), .B0(N67), .B1(n50), .Y(n165) );
  AOI22X1 U91 ( .A0(N98), .A1(n57), .B0(N66), .B1(n50), .Y(n171) );
  AOI22X1 U92 ( .A0(N97), .A1(n57), .B0(N65), .B1(n50), .Y(n177) );
  AOI22X1 U93 ( .A0(N96), .A1(n57), .B0(N64), .B1(n50), .Y(n189) );
  AOI22X1 U94 ( .A0(N95), .A1(n57), .B0(N63), .B1(n50), .Y(n195) );
  AOI22X1 U95 ( .A0(N94), .A1(n57), .B0(N62), .B1(n50), .Y(n201) );
  AOI22X1 U96 ( .A0(N93), .A1(n57), .B0(N61), .B1(n50), .Y(n207) );
  AOI22X1 U97 ( .A0(N92), .A1(n52), .B0(N60), .B1(n50), .Y(n213) );
  AOI2BB2X1 U98 ( .B0(N214), .B1(n44), .A0N(n48), .A1N(n297), .Y(n70) );
  AOI2BB2X1 U99 ( .B0(N212), .B1(n44), .A0N(n47), .A1N(n299), .Y(n82) );
  AOI221XL U100 ( .A0(N86), .A1(n52), .B0(N54), .B1(n58), .C0(n59), .Y(n56) );
  OAI2BB2XL U101 ( .B0(n296), .B1(n46), .A0N(N215), .A1N(n61), .Y(n59) );
  AOI22X1 U102 ( .A0(N91), .A1(n52), .B0(N59), .B1(n50), .Y(n219) );
  AOI22X1 U103 ( .A0(N85), .A1(n51), .B0(N53), .B1(n49), .Y(n69) );
  AOI22X1 U104 ( .A0(N84), .A1(n51), .B0(N52), .B1(n49), .Y(n75) );
  AOI22X1 U105 ( .A0(N90), .A1(n52), .B0(N58), .B1(n58), .Y(n225) );
  AOI22X1 U106 ( .A0(N89), .A1(n52), .B0(N57), .B1(n58), .Y(n231) );
  AOI22X1 U107 ( .A0(N88), .A1(n52), .B0(N56), .B1(n58), .Y(n237) );
  AOI22X1 U108 ( .A0(N87), .A1(n52), .B0(N55), .B1(n58), .Y(n243) );
  AOI2BB2X1 U109 ( .B0(N236), .B1(n45), .A0N(n48), .A1N(n275), .Y(n112) );
  AOI2BB2X1 U110 ( .B0(N235), .B1(n44), .A0N(n48), .A1N(n276), .Y(n124) );
  AOI2BB2X1 U111 ( .B0(N234), .B1(n44), .A0N(n48), .A1N(n277), .Y(n130) );
  AOI2BB2X1 U112 ( .B0(N233), .B1(n44), .A0N(n48), .A1N(n278), .Y(n136) );
  AOI2BB2X1 U113 ( .B0(N232), .B1(n44), .A0N(n48), .A1N(n279), .Y(n142) );
  AOI2BB2X1 U114 ( .B0(N231), .B1(n45), .A0N(n48), .A1N(n280), .Y(n148) );
  AOI2BB2X1 U115 ( .B0(N230), .B1(n45), .A0N(n48), .A1N(n281), .Y(n154) );
  AOI2BB2X1 U116 ( .B0(N229), .B1(n45), .A0N(n48), .A1N(n282), .Y(n160) );
  AOI2BB2X1 U117 ( .B0(N228), .B1(n45), .A0N(n48), .A1N(n283), .Y(n166) );
  AOI2BB2X1 U118 ( .B0(N227), .B1(n45), .A0N(n48), .A1N(n284), .Y(n172) );
  AOI2BB2X1 U119 ( .B0(N226), .B1(n45), .A0N(n48), .A1N(n285), .Y(n178) );
  AOI2BB2X1 U120 ( .B0(N224), .B1(n45), .A0N(n48), .A1N(n287), .Y(n196) );
  AOI2BB2X1 U121 ( .B0(N223), .B1(n45), .A0N(n48), .A1N(n288), .Y(n202) );
  AOI2BB2X1 U122 ( .B0(N222), .B1(n45), .A0N(n48), .A1N(n289), .Y(n208) );
  AOI2BB2X1 U123 ( .B0(N213), .B1(n44), .A0N(n47), .A1N(n298), .Y(n76) );
  AOI2BB2X1 U124 ( .B0(N237), .B1(n44), .A0N(n47), .A1N(n274), .Y(n106) );
  AOI2BB2X1 U125 ( .B0(N221), .B1(n61), .A0N(n48), .A1N(n290), .Y(n214) );
  AOI2BB2X1 U126 ( .B0(N220), .B1(n61), .A0N(n48), .A1N(n291), .Y(n220) );
  AOI2BB2X1 U127 ( .B0(N219), .B1(n61), .A0N(n60), .A1N(n292), .Y(n226) );
  AOI2BB2X1 U128 ( .B0(N218), .B1(n44), .A0N(n48), .A1N(n293), .Y(n232) );
  AOI2BB2X1 U129 ( .B0(N217), .B1(n61), .A0N(n60), .A1N(n294), .Y(n238) );
  AOI2BB2X1 U130 ( .B0(N216), .B1(n61), .A0N(n60), .A1N(n295), .Y(n244) );
  AOI2BB2X1 U131 ( .B0(N225), .B1(n45), .A0N(n48), .A1N(n286), .Y(n190) );
  CLKINVX1 U132 ( .A(ctrl[1]), .Y(n300) );
  NOR2BX1 U133 ( .AN(ctrl[2]), .B(ctrl[3]), .Y(n253) );
  CLKINVX1 U134 ( .A(ctrl[0]), .Y(n301) );
  NOR2X1 U135 ( .A(ctrl[3]), .B(ctrl[2]), .Y(n254) );
  NAND3X1 U136 ( .A(ctrl[0]), .B(n254), .C(ctrl[1]), .Y(n64) );
  AND3X2 U137 ( .A(n253), .B(n300), .C(ctrl[0]), .Y(n61) );
  AND3X2 U138 ( .A(n254), .B(n301), .C(ctrl[1]), .Y(n58) );
  AND3X2 U139 ( .A(n253), .B(n301), .C(ctrl[1]), .Y(n57) );
  NOR3BXL U140 ( .AN(ctrl[3]), .B(ctrl[1]), .C(ctrl[2]), .Y(n258) );
  NAND3X1 U141 ( .A(n254), .B(n300), .C(ctrl[0]), .Y(n60) );
  AND2X2 U142 ( .A(n258), .B(ctrl[0]), .Y(n67) );
  AOI22X1 U143 ( .A0(N83), .A1(n51), .B0(N51), .B1(n49), .Y(n81) );
  AOI22X1 U144 ( .A0(N108), .A1(n51), .B0(N76), .B1(n49), .Y(n105) );
  INVX3 U145 ( .A(n265), .Y(n264) );
  AOI2BB2X1 U146 ( .B0(N211), .B1(n44), .A0N(n46), .A1N(n259), .Y(n88) );
  AOI2BB2X1 U147 ( .B0(N210), .B1(n44), .A0N(n46), .A1N(n261), .Y(n94) );
  OAI2BB2XL U148 ( .B0(n46), .B1(n269), .A0N(N206), .A1N(n61), .Y(n252) );
  AOI221XL U149 ( .A0(n270), .A1(n255), .B0(n256), .B1(n271), .C0(n257), .Y(
        n250) );
  OAI22XL U150 ( .A0(n41), .A1(n269), .B0(n268), .B1(n39), .Y(n256) );
  OAI221XL U151 ( .A0(n268), .A1(n41), .B0(n37), .B1(n269), .C0(n46), .Y(n255)
         );
  AND4X1 U152 ( .A(N205), .B(ctrl[1]), .C(ctrl[0]), .D(n253), .Y(n257) );
  AOI2BB2X1 U153 ( .B0(N209), .B1(n44), .A0N(n48), .A1N(n263), .Y(n100) );
  AOI2BB2X1 U154 ( .B0(N208), .B1(n44), .A0N(n48), .A1N(n265), .Y(n118) );
  AOI2BB2X1 U155 ( .B0(N207), .B1(n45), .A0N(n47), .A1N(n267), .Y(n184) );
  OAI221XL U156 ( .A0(n31), .A1(n42), .B0(n37), .B1(n275), .C0(n46), .Y(n115)
         );
  OAI221XL U157 ( .A0(n30), .A1(n42), .B0(n37), .B1(n276), .C0(n46), .Y(n127)
         );
  OAI221XL U158 ( .A0(n29), .A1(n42), .B0(n37), .B1(n277), .C0(n46), .Y(n133)
         );
  OAI221XL U159 ( .A0(n28), .A1(n42), .B0(n37), .B1(n278), .C0(n47), .Y(n139)
         );
  OAI221XL U160 ( .A0(n27), .A1(n42), .B0(n38), .B1(n279), .C0(n46), .Y(n145)
         );
  OAI221XL U161 ( .A0(n26), .A1(n42), .B0(n38), .B1(n280), .C0(n46), .Y(n151)
         );
  OAI221XL U162 ( .A0(n25), .A1(n42), .B0(n38), .B1(n281), .C0(n47), .Y(n157)
         );
  OAI221XL U163 ( .A0(n24), .A1(n42), .B0(n38), .B1(n282), .C0(n47), .Y(n163)
         );
  OAI221XL U164 ( .A0(n23), .A1(n42), .B0(n38), .B1(n283), .C0(n47), .Y(n169)
         );
  OAI221XL U165 ( .A0(n22), .A1(n42), .B0(n38), .B1(n284), .C0(n47), .Y(n175)
         );
  OAI221XL U166 ( .A0(n21), .A1(n42), .B0(n38), .B1(n285), .C0(n47), .Y(n181)
         );
  OAI221XL U167 ( .A0(n20), .A1(n42), .B0(n38), .B1(n286), .C0(n47), .Y(n193)
         );
  OAI221XL U168 ( .A0(n19), .A1(n41), .B0(n38), .B1(n287), .C0(n47), .Y(n199)
         );
  OAI221XL U169 ( .A0(n12), .A1(n41), .B0(n38), .B1(n288), .C0(n47), .Y(n205)
         );
  OAI221XL U170 ( .A0(n11), .A1(n41), .B0(n38), .B1(n289), .C0(n47), .Y(n211)
         );
  OAI221XL U171 ( .A0(n10), .A1(n41), .B0(n38), .B1(n290), .C0(n47), .Y(n217)
         );
  OAI221XL U172 ( .A0(n4), .A1(n41), .B0(n296), .B1(n37), .C0(n46), .Y(n62) );
  OAI221XL U173 ( .A0(n9), .A1(n41), .B0(n66), .B1(n291), .C0(n47), .Y(n223)
         );
  OAI221XL U174 ( .A0(n8), .A1(n41), .B0(n66), .B1(n292), .C0(n47), .Y(n229)
         );
  OAI221XL U175 ( .A0(n7), .A1(n41), .B0(n38), .B1(n293), .C0(n47), .Y(n235)
         );
  OAI221XL U176 ( .A0(n6), .A1(n41), .B0(n38), .B1(n294), .C0(n47), .Y(n241)
         );
  OAI221XL U177 ( .A0(n5), .A1(n41), .B0(n37), .B1(n295), .C0(n47), .Y(n247)
         );
  OAI221XL U178 ( .A0(n3), .A1(n41), .B0(n37), .B1(n297), .C0(n46), .Y(n73) );
  OAI221XL U179 ( .A0(n2), .A1(n41), .B0(n37), .B1(n298), .C0(n46), .Y(n79) );
  OAI221XL U180 ( .A0(n1), .A1(n41), .B0(n37), .B1(n299), .C0(n46), .Y(n85) );
  OAI221XL U181 ( .A0(n53), .A1(n41), .B0(n37), .B1(n259), .C0(n46), .Y(n91)
         );
  OAI221XL U182 ( .A0(n260), .A1(n42), .B0(n37), .B1(n261), .C0(n46), .Y(n97)
         );
  OAI221XL U183 ( .A0(n262), .A1(n42), .B0(n37), .B1(n263), .C0(n46), .Y(n103)
         );
  OAI221XL U184 ( .A0(n264), .A1(n43), .B0(n37), .B1(n265), .C0(n46), .Y(n121)
         );
  OAI221XL U185 ( .A0(n32), .A1(n42), .B0(n37), .B1(n274), .C0(n46), .Y(n109)
         );
  AOI2BB2X1 U186 ( .B0(y[1]), .B1(n187), .A0N(n188), .A1N(y[1]), .Y(n186) );
  OA22X1 U187 ( .A0(n42), .A1(n267), .B0(n266), .B1(n39), .Y(n188) );
  OAI221XL U188 ( .A0(n266), .A1(n42), .B0(n38), .B1(n267), .C0(n47), .Y(n187)
         );
  CLKINVX1 U189 ( .A(n4), .Y(n296) );
  CLKINVX1 U190 ( .A(n19), .Y(n287) );
  CLKINVX1 U191 ( .A(n31), .Y(n275) );
  CLKINVX1 U192 ( .A(n27), .Y(n279) );
  CLKINVX1 U193 ( .A(n25), .Y(n281) );
  CLKINVX1 U194 ( .A(n9), .Y(n291) );
  CLKINVX1 U195 ( .A(n11), .Y(n289) );
  CLKINVX1 U196 ( .A(n12), .Y(n288) );
  CLKINVX1 U197 ( .A(n28), .Y(n278) );
  CLKINVX1 U198 ( .A(n26), .Y(n280) );
  CLKINVX1 U199 ( .A(n24), .Y(n282) );
  CLKINVX1 U200 ( .A(n23), .Y(n283) );
  CLKINVX1 U201 ( .A(n10), .Y(n290) );
  CLKINVX1 U202 ( .A(n2), .Y(n298) );
  CLKINVX1 U203 ( .A(n21), .Y(n285) );
  CLKINVX1 U204 ( .A(n1), .Y(n299) );
  CLKINVX1 U205 ( .A(n32), .Y(n274) );
  CLKINVX1 U206 ( .A(n22), .Y(n284) );
  CLKINVX1 U207 ( .A(n20), .Y(n286) );
  CLKINVX1 U208 ( .A(n3), .Y(n297) );
  CLKINVX1 U209 ( .A(n30), .Y(n276) );
  CLKINVX1 U210 ( .A(n29), .Y(n277) );
  CLKINVX1 U211 ( .A(n8), .Y(n292) );
  CLKINVX1 U212 ( .A(n7), .Y(n293) );
  CLKINVX1 U213 ( .A(n6), .Y(n294) );
  CLKINVX1 U214 ( .A(n5), .Y(n295) );
  OA22X1 U215 ( .A0(n43), .A1(n259), .B0(n53), .B1(n40), .Y(n92) );
  OA22X1 U216 ( .A0(n43), .A1(n261), .B0(n260), .B1(n40), .Y(n98) );
  OA22X1 U217 ( .A0(n43), .A1(n263), .B0(n262), .B1(n40), .Y(n104) );
  OA22X1 U218 ( .A0(n43), .A1(n265), .B0(n264), .B1(n40), .Y(n122) );
  OA22X1 U219 ( .A0(n43), .A1(n275), .B0(n31), .B1(n40), .Y(n116) );
  OA22X1 U220 ( .A0(n43), .A1(n278), .B0(n28), .B1(n40), .Y(n140) );
  OA22X1 U221 ( .A0(n43), .A1(n279), .B0(n27), .B1(n40), .Y(n146) );
  OA22X1 U222 ( .A0(n41), .A1(n284), .B0(n22), .B1(n39), .Y(n176) );
  OA22X1 U223 ( .A0(n41), .A1(n287), .B0(n19), .B1(n39), .Y(n200) );
  OA22X1 U224 ( .A0(n43), .A1(n276), .B0(n30), .B1(n40), .Y(n128) );
  OA22X1 U225 ( .A0(n43), .A1(n277), .B0(n29), .B1(n40), .Y(n134) );
  OA22X1 U226 ( .A0(n43), .A1(n280), .B0(n26), .B1(n39), .Y(n152) );
  OA22X1 U227 ( .A0(n43), .A1(n281), .B0(n25), .B1(n39), .Y(n158) );
  OA22X1 U228 ( .A0(n43), .A1(n282), .B0(n24), .B1(n39), .Y(n164) );
  OA22X1 U229 ( .A0(n41), .A1(n283), .B0(n23), .B1(n39), .Y(n170) );
  OA22X1 U230 ( .A0(n43), .A1(n285), .B0(n21), .B1(n39), .Y(n182) );
  OA22X1 U231 ( .A0(n42), .A1(n286), .B0(n20), .B1(n39), .Y(n194) );
  OA22X1 U232 ( .A0(n64), .A1(n288), .B0(n12), .B1(n39), .Y(n206) );
  OA22X1 U233 ( .A0(n41), .A1(n289), .B0(n11), .B1(n39), .Y(n212) );
  OA22X1 U234 ( .A0(n42), .A1(n290), .B0(n10), .B1(n39), .Y(n218) );
  OA22X1 U235 ( .A0(n43), .A1(n291), .B0(n9), .B1(n39), .Y(n224) );
  OA22X1 U236 ( .A0(n42), .A1(n292), .B0(n8), .B1(n39), .Y(n230) );
  OA22X1 U237 ( .A0(n42), .A1(n293), .B0(n7), .B1(n39), .Y(n236) );
  OA22X1 U238 ( .A0(n41), .A1(n294), .B0(n6), .B1(n39), .Y(n242) );
  OA22X1 U239 ( .A0(n43), .A1(n295), .B0(n5), .B1(n39), .Y(n248) );
  OA22X1 U240 ( .A0(n43), .A1(n296), .B0(n4), .B1(n40), .Y(n63) );
  OA22X1 U241 ( .A0(n43), .A1(n297), .B0(n3), .B1(n40), .Y(n74) );
  OA22X1 U242 ( .A0(n43), .A1(n298), .B0(n2), .B1(n40), .Y(n80) );
  OA22X1 U243 ( .A0(n43), .A1(n299), .B0(n1), .B1(n40), .Y(n86) );
  OA22X1 U244 ( .A0(n43), .A1(n274), .B0(n32), .B1(n40), .Y(n110) );
  NAND4X1 U245 ( .A(n105), .B(n106), .C(n107), .D(n108), .Y(out[31]) );
  AOI2BB2X1 U246 ( .B0(y[31]), .B1(n109), .A0N(n110), .A1N(y[31]), .Y(n108) );
  NAND4X1 U247 ( .A(n111), .B(n112), .C(n113), .D(n114), .Y(out[30]) );
  AOI2BB2X1 U248 ( .B0(y[30]), .B1(n115), .A0N(n116), .A1N(y[30]), .Y(n114) );
  NAND4X1 U249 ( .A(n129), .B(n130), .C(n131), .D(n132), .Y(out[28]) );
  AOI2BB2X1 U250 ( .B0(y[28]), .B1(n133), .A0N(n134), .A1N(y[28]), .Y(n132) );
  NAND4X1 U251 ( .A(n141), .B(n142), .C(n143), .D(n144), .Y(out[26]) );
  AOI2BB2X1 U252 ( .B0(y[26]), .B1(n145), .A0N(n146), .A1N(y[26]), .Y(n144) );
  NAND4X1 U253 ( .A(n153), .B(n154), .C(n155), .D(n156), .Y(out[24]) );
  AOI2BB2X1 U254 ( .B0(y[24]), .B1(n157), .A0N(n158), .A1N(y[24]), .Y(n156) );
  NAND4X1 U255 ( .A(n135), .B(n136), .C(n137), .D(n138), .Y(out[27]) );
  AOI2BB2X1 U256 ( .B0(y[27]), .B1(n139), .A0N(n140), .A1N(y[27]), .Y(n138) );
  NAND4X1 U257 ( .A(n147), .B(n148), .C(n149), .D(n150), .Y(out[25]) );
  AOI2BB2X1 U258 ( .B0(y[25]), .B1(n151), .A0N(n152), .A1N(y[25]), .Y(n150) );
  NAND4X1 U259 ( .A(n123), .B(n124), .C(n125), .D(n126), .Y(out[29]) );
  AOI2BB2X1 U260 ( .B0(y[29]), .B1(n127), .A0N(n128), .A1N(y[29]), .Y(n126) );
  CLKBUFX3 U261 ( .A(x[6]), .Y(n1) );
  NAND4X1 U262 ( .A(n159), .B(n160), .C(n161), .D(n162), .Y(out[23]) );
  AOI2BB2X1 U263 ( .B0(y[23]), .B1(n163), .A0N(n164), .A1N(y[23]), .Y(n162) );
  NAND4X1 U264 ( .A(n165), .B(n166), .C(n167), .D(n168), .Y(out[22]) );
  AOI2BB2X1 U265 ( .B0(y[22]), .B1(n169), .A0N(n170), .A1N(y[22]), .Y(n168) );
  NAND4X1 U266 ( .A(n177), .B(n178), .C(n179), .D(n180), .Y(out[20]) );
  AOI2BB2X1 U267 ( .B0(y[20]), .B1(n181), .A0N(n182), .A1N(y[20]), .Y(n180) );
  NAND4X1 U268 ( .A(n189), .B(n190), .C(n191), .D(n192), .Y(out[19]) );
  AOI2BB2X1 U269 ( .B0(y[19]), .B1(n193), .A0N(n194), .A1N(y[19]), .Y(n192) );
  NAND4X1 U270 ( .A(n201), .B(n202), .C(n203), .D(n204), .Y(out[17]) );
  AOI2BB2X1 U271 ( .B0(y[17]), .B1(n205), .A0N(n206), .A1N(y[17]), .Y(n204) );
  NAND4X1 U272 ( .A(n207), .B(n208), .C(n209), .D(n210), .Y(out[16]) );
  AOI2BB2X1 U273 ( .B0(y[16]), .B1(n211), .A0N(n212), .A1N(y[16]), .Y(n210) );
  CLKBUFX3 U274 ( .A(x[9]), .Y(n4) );
  CLKBUFX3 U275 ( .A(x[7]), .Y(n2) );
  CLKBUFX3 U276 ( .A(x[14]), .Y(n9) );
  CLKBUFX3 U277 ( .A(x[8]), .Y(n3) );
  CLKBUFX3 U278 ( .A(x[12]), .Y(n7) );
  CLKBUFX3 U279 ( .A(x[11]), .Y(n6) );
  CLKBUFX3 U280 ( .A(x[13]), .Y(n8) );
  CLKBUFX3 U281 ( .A(x[10]), .Y(n5) );
  NAND4X1 U282 ( .A(n213), .B(n214), .C(n215), .D(n216), .Y(out[15]) );
  AOI2BB2X1 U283 ( .B0(y[15]), .B1(n217), .A0N(n218), .A1N(y[15]), .Y(n216) );
  NAND4X1 U284 ( .A(n171), .B(n172), .C(n173), .D(n174), .Y(out[21]) );
  AOI2BB2X1 U285 ( .B0(y[21]), .B1(n175), .A0N(n176), .A1N(y[21]), .Y(n174) );
  NAND4X1 U286 ( .A(n195), .B(n196), .C(n197), .D(n198), .Y(out[18]) );
  AOI2BB2X1 U287 ( .B0(y[18]), .B1(n199), .A0N(n200), .A1N(y[18]), .Y(n198) );
  CLKBUFX3 U288 ( .A(x[24]), .Y(n25) );
  NAND4X1 U289 ( .A(n219), .B(n220), .C(n221), .D(n222), .Y(out[14]) );
  AOI2BB2X1 U290 ( .B0(y[14]), .B1(n223), .A0N(n224), .A1N(y[14]), .Y(n222) );
  NAND4X1 U291 ( .A(n225), .B(n226), .C(n227), .D(n228), .Y(out[13]) );
  AOI2BB2X1 U292 ( .B0(y[13]), .B1(n229), .A0N(n230), .A1N(y[13]), .Y(n228) );
  NAND4X1 U293 ( .A(n237), .B(n238), .C(n239), .D(n240), .Y(out[11]) );
  AOI2BB2X1 U294 ( .B0(y[11]), .B1(n241), .A0N(n242), .A1N(y[11]), .Y(n240) );
  NAND4X1 U295 ( .A(n243), .B(n244), .C(n245), .D(n246), .Y(out[10]) );
  AOI2BB2X1 U296 ( .B0(y[10]), .B1(n247), .A0N(n248), .A1N(y[10]), .Y(n246) );
  NAND4X1 U297 ( .A(n69), .B(n70), .C(n71), .D(n72), .Y(out[8]) );
  AOI2BB2X1 U298 ( .B0(y[8]), .B1(n73), .A0N(n74), .A1N(y[8]), .Y(n72) );
  NAND4X1 U299 ( .A(n81), .B(n82), .C(n83), .D(n84), .Y(out[6]) );
  AOI2BB2X1 U300 ( .B0(y[6]), .B1(n85), .A0N(n86), .A1N(y[6]), .Y(n84) );
  NAND4X1 U301 ( .A(n87), .B(n88), .C(n89), .D(n90), .Y(out[5]) );
  AOI2BB2X1 U302 ( .B0(n273), .B1(n91), .A0N(n92), .A1N(n273), .Y(n90) );
  NAND4X1 U303 ( .A(n99), .B(n100), .C(n101), .D(n102), .Y(out[3]) );
  AOI2BB2X1 U304 ( .B0(y[3]), .B1(n103), .A0N(n104), .A1N(y[3]), .Y(n102) );
  NAND4X1 U305 ( .A(n117), .B(n118), .C(n119), .D(n120), .Y(out[2]) );
  AOI2BB2X1 U306 ( .B0(y[2]), .B1(n121), .A0N(n122), .A1N(y[2]), .Y(n120) );
  CLKBUFX3 U307 ( .A(x[17]), .Y(n12) );
  CLKBUFX3 U308 ( .A(x[18]), .Y(n19) );
  CLKBUFX3 U309 ( .A(x[23]), .Y(n24) );
  CLKBUFX3 U310 ( .A(x[15]), .Y(n10) );
  CLKBUFX3 U311 ( .A(x[16]), .Y(n11) );
  CLKBUFX3 U312 ( .A(x[31]), .Y(n32) );
  NAND4X1 U313 ( .A(n183), .B(n184), .C(n185), .D(n186), .Y(out[1]) );
  AOI22X1 U314 ( .A0(N78), .A1(n57), .B0(N46), .B1(n50), .Y(n183) );
  NAND4X1 U315 ( .A(n75), .B(n76), .C(n77), .D(n78), .Y(out[7]) );
  AOI2BB2X1 U316 ( .B0(y[7]), .B1(n79), .A0N(n80), .A1N(y[7]), .Y(n78) );
  NAND4X1 U317 ( .A(n231), .B(n232), .C(n233), .D(n234), .Y(out[12]) );
  AOI2BB2X1 U318 ( .B0(y[12]), .B1(n235), .A0N(n236), .A1N(y[12]), .Y(n234) );
  NAND3X1 U319 ( .A(n249), .B(n250), .C(n251), .Y(out[0]) );
  AOI221XL U320 ( .A0(N77), .A1(n52), .B0(N45), .B1(n58), .C0(n252), .Y(n251)
         );
  CLKBUFX3 U321 ( .A(x[30]), .Y(n31) );
  CLKBUFX3 U322 ( .A(x[26]), .Y(n27) );
  CLKBUFX3 U323 ( .A(x[25]), .Y(n26) );
  CLKBUFX3 U324 ( .A(x[27]), .Y(n28) );
  CLKBUFX3 U325 ( .A(x[22]), .Y(n23) );
  CLKBUFX3 U326 ( .A(x[20]), .Y(n21) );
  CLKBUFX3 U327 ( .A(x[21]), .Y(n22) );
  CLKBUFX3 U328 ( .A(x[19]), .Y(n20) );
  CLKBUFX3 U329 ( .A(x[28]), .Y(n29) );
  CLKBUFX3 U330 ( .A(x[29]), .Y(n30) );
  NAND4X1 U331 ( .A(n93), .B(n94), .C(n95), .D(n96), .Y(out[4]) );
  AOI2BB2X1 U332 ( .B0(n272), .B1(n97), .A0N(n98), .A1N(n272), .Y(n96) );
  NAND3X1 U333 ( .A(n54), .B(n55), .C(n56), .Y(out[9]) );
  AOI2BB2X1 U334 ( .B0(y[9]), .B1(n62), .A0N(n63), .A1N(y[9]), .Y(n55) );
endmodule


module mul_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [32:1] carry;

  ADDFXL U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDFXL U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(SUM[32]), .S(
        SUM[31]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFXL U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module mul_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [33:0] carry;

  ADDFXL U2_31 ( .A(A[31]), .B(n9), .CI(carry[31]), .CO(carry[32]), .S(
        DIFF[31]) );
  ADDFXL U2_30 ( .A(A[30]), .B(n8), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  ADDFXL U2_29 ( .A(A[29]), .B(n7), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  ADDFXL U2_28 ( .A(A[28]), .B(n6), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  ADDFXL U2_27 ( .A(A[27]), .B(n5), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  ADDFXL U2_26 ( .A(A[26]), .B(n4), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  ADDFXL U2_25 ( .A(A[25]), .B(n3), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  ADDFXL U2_24 ( .A(A[24]), .B(n33), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  ADDFXL U2_23 ( .A(A[23]), .B(n32), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  ADDFXL U2_22 ( .A(A[22]), .B(n31), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  ADDFXL U2_21 ( .A(A[21]), .B(n30), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  ADDFXL U2_20 ( .A(A[20]), .B(n29), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  ADDFXL U2_19 ( .A(A[19]), .B(n28), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  ADDFXL U2_18 ( .A(A[18]), .B(n27), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  ADDFXL U2_17 ( .A(A[17]), .B(n26), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  ADDFXL U2_16 ( .A(A[16]), .B(n25), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  ADDFXL U2_15 ( .A(A[15]), .B(n24), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n23), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n22), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n21), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n20), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n19), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n18), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n17), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  ADDFXL U2_7 ( .A(A[7]), .B(n16), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n15), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n14), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n12), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n11), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n10), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  CLKINVX1 U1 ( .A(B[0]), .Y(n2) );
  CLKINVX1 U2 ( .A(B[1]), .Y(n10) );
  NAND2X1 U3 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U4 ( .A(A[0]), .Y(n1) );
  CLKINVX1 U5 ( .A(B[2]), .Y(n11) );
  CLKINVX1 U6 ( .A(B[3]), .Y(n12) );
  CLKINVX1 U7 ( .A(B[4]), .Y(n13) );
  CLKINVX1 U8 ( .A(B[5]), .Y(n14) );
  CLKINVX1 U9 ( .A(B[6]), .Y(n15) );
  CLKINVX1 U10 ( .A(B[7]), .Y(n16) );
  CLKINVX1 U11 ( .A(B[8]), .Y(n17) );
  CLKINVX1 U12 ( .A(B[9]), .Y(n18) );
  CLKINVX1 U13 ( .A(B[10]), .Y(n19) );
  CLKINVX1 U14 ( .A(B[11]), .Y(n20) );
  CLKINVX1 U15 ( .A(B[12]), .Y(n21) );
  CLKINVX1 U16 ( .A(B[13]), .Y(n22) );
  CLKINVX1 U17 ( .A(B[14]), .Y(n23) );
  CLKINVX1 U18 ( .A(B[15]), .Y(n24) );
  CLKINVX1 U19 ( .A(B[16]), .Y(n25) );
  CLKINVX1 U20 ( .A(B[17]), .Y(n26) );
  CLKINVX1 U21 ( .A(B[18]), .Y(n27) );
  CLKINVX1 U22 ( .A(B[19]), .Y(n28) );
  CLKINVX1 U23 ( .A(B[20]), .Y(n29) );
  CLKINVX1 U24 ( .A(B[21]), .Y(n30) );
  CLKINVX1 U25 ( .A(B[22]), .Y(n31) );
  CLKINVX1 U26 ( .A(B[23]), .Y(n32) );
  CLKINVX1 U27 ( .A(B[24]), .Y(n33) );
  CLKINVX1 U28 ( .A(B[25]), .Y(n3) );
  CLKINVX1 U29 ( .A(B[26]), .Y(n4) );
  CLKINVX1 U30 ( .A(B[27]), .Y(n5) );
  CLKINVX1 U31 ( .A(B[28]), .Y(n6) );
  CLKINVX1 U32 ( .A(B[29]), .Y(n7) );
  CLKINVX1 U33 ( .A(B[30]), .Y(n8) );
  CLKINVX1 U34 ( .A(B[31]), .Y(n9) );
  XNOR2X1 U35 ( .A(n2), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U36 ( .A(carry[32]), .Y(DIFF[32]) );
endmodule


module mul ( clk, rst, mul, multiplicand, LO, next_HI, next_LO, mul_stall );
  input [31:0] multiplicand;
  input [31:0] LO;
  output [31:0] next_HI;
  output [31:0] next_LO;
  input clk, rst, mul;
  output mul_stall;
  wire   n37, state_w, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87,
         N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N107,
         N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118,
         N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129,
         N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N173,
         N174, N175, N176, N177, N178, state_r, n7, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, \add_56/carry[5] ,
         \add_56/carry[4] , \add_56/carry[3] , \add_56/carry[2] , n3, n4, n5,
         n6, n8, n22, n23, n24, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36;
  wire   [5:0] mul_iter_r;
  wire   [31:0] HI_w;
  wire   [31:0] LO_w;

  mul_DW01_add_0 add_49 ( .A({1'b0, next_HI}), .B({1'b0, N41, N40, N39, N38, 
        N37, N36, N35, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, 
        N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75}), 
        .CI(1'b0), .SUM({N139, N138, N137, N136, N135, N134, N133, N132, N131, 
        N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, 
        N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107}) );
  mul_DW01_sub_0 sub_45 ( .A({1'b0, next_HI}), .B({1'b0, N41, N40, N39, N38, 
        N37, N36, N35, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, 
        N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75}), 
        .CI(1'b0), .DIFF({N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, 
        N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, 
        N50, N49, N48, N47, N46, N45, N44, N43, N42}) );
  ADDHXL \add_56/U1_1_4  ( .A(mul_iter_r[4]), .B(\add_56/carry[4] ), .CO(
        \add_56/carry[5] ), .S(N177) );
  ADDHXL \add_56/U1_1_1  ( .A(mul_iter_r[1]), .B(mul_iter_r[0]), .CO(
        \add_56/carry[2] ), .S(N174) );
  ADDHXL \add_56/U1_1_3  ( .A(mul_iter_r[3]), .B(\add_56/carry[3] ), .CO(
        \add_56/carry[4] ), .S(N176) );
  ADDHXL \add_56/U1_1_2  ( .A(mul_iter_r[2]), .B(\add_56/carry[2] ), .CO(
        \add_56/carry[3] ), .S(N175) );
  DFFSX1 \mul_iter_r_reg[5]  ( .D(n20), .CK(clk), .SN(n33), .Q(mul_iter_r[5]), 
        .QN(n7) );
  DFFRX1 state_r_reg ( .D(state_w), .CK(clk), .RN(n28), .Q(state_r) );
  DFFRX1 \mul_iter_r_reg[4]  ( .D(n19), .CK(clk), .RN(n28), .Q(mul_iter_r[4])
         );
  DFFRX1 \mul_iter_r_reg[3]  ( .D(n18), .CK(clk), .RN(n28), .Q(mul_iter_r[3])
         );
  DFFRX1 \mul_iter_r_reg[2]  ( .D(n17), .CK(clk), .RN(n28), .Q(mul_iter_r[2])
         );
  DFFRX1 \mul_iter_r_reg[1]  ( .D(n16), .CK(clk), .RN(n28), .Q(mul_iter_r[1])
         );
  DFFRX1 \mul_iter_r_reg[0]  ( .D(n21), .CK(clk), .RN(n28), .Q(mul_iter_r[0]), 
        .QN(N173) );
  DFFRX1 \LO_r_reg[16]  ( .D(LO_w[16]), .CK(clk), .RN(n29), .Q(next_LO[16]) );
  DFFRX1 \LO_r_reg[15]  ( .D(LO_w[15]), .CK(clk), .RN(n30), .Q(next_LO[15]) );
  DFFRX1 \LO_r_reg[14]  ( .D(LO_w[14]), .CK(clk), .RN(n30), .Q(next_LO[14]) );
  DFFRX1 \LO_r_reg[13]  ( .D(LO_w[13]), .CK(clk), .RN(n30), .Q(next_LO[13]) );
  DFFRX1 \LO_r_reg[12]  ( .D(LO_w[12]), .CK(clk), .RN(n30), .Q(next_LO[12]) );
  DFFRX1 \LO_r_reg[11]  ( .D(LO_w[11]), .CK(clk), .RN(n30), .Q(next_LO[11]) );
  DFFRX1 \LO_r_reg[10]  ( .D(LO_w[10]), .CK(clk), .RN(n30), .Q(next_LO[10]) );
  DFFRX1 \LO_r_reg[0]  ( .D(LO_w[0]), .CK(clk), .RN(n28), .Q(n37) );
  DFFRX1 \LO_r_reg[9]  ( .D(LO_w[9]), .CK(clk), .RN(n30), .Q(next_LO[9]) );
  DFFRX1 \LO_r_reg[30]  ( .D(LO_w[30]), .CK(clk), .RN(n28), .Q(next_LO[30]) );
  DFFRX1 \LO_r_reg[29]  ( .D(LO_w[29]), .CK(clk), .RN(n28), .Q(next_LO[29]) );
  DFFRX1 \LO_r_reg[28]  ( .D(LO_w[28]), .CK(clk), .RN(n28), .Q(next_LO[28]) );
  DFFRX1 \LO_r_reg[2]  ( .D(LO_w[2]), .CK(clk), .RN(n31), .Q(next_LO[2]) );
  DFFRX1 \LO_r_reg[8]  ( .D(LO_w[8]), .CK(clk), .RN(n30), .Q(next_LO[8]) );
  DFFRX1 \LO_r_reg[7]  ( .D(LO_w[7]), .CK(clk), .RN(n30), .Q(next_LO[7]) );
  DFFRX1 \LO_r_reg[6]  ( .D(LO_w[6]), .CK(clk), .RN(n30), .Q(next_LO[6]) );
  DFFRX1 \LO_r_reg[5]  ( .D(LO_w[5]), .CK(clk), .RN(n30), .Q(next_LO[5]) );
  DFFRX1 \LO_r_reg[4]  ( .D(LO_w[4]), .CK(clk), .RN(n30), .Q(next_LO[4]) );
  DFFRX1 \LO_r_reg[3]  ( .D(LO_w[3]), .CK(clk), .RN(n31), .Q(next_LO[3]) );
  DFFRX1 \LO_r_reg[19]  ( .D(LO_w[19]), .CK(clk), .RN(n29), .Q(next_LO[19]) );
  DFFRX1 \LO_r_reg[18]  ( .D(LO_w[18]), .CK(clk), .RN(n29), .Q(next_LO[18]) );
  DFFRX1 \LO_r_reg[17]  ( .D(LO_w[17]), .CK(clk), .RN(n29), .Q(next_LO[17]) );
  DFFRX1 \LO_r_reg[1]  ( .D(LO_w[1]), .CK(clk), .RN(n31), .Q(next_LO[1]) );
  DFFRX1 \LO_r_reg[27]  ( .D(LO_w[27]), .CK(clk), .RN(n29), .Q(next_LO[27]) );
  DFFRX1 \LO_r_reg[26]  ( .D(LO_w[26]), .CK(clk), .RN(n29), .Q(next_LO[26]) );
  DFFRX1 \LO_r_reg[25]  ( .D(LO_w[25]), .CK(clk), .RN(n29), .Q(next_LO[25]) );
  DFFRX1 \LO_r_reg[24]  ( .D(LO_w[24]), .CK(clk), .RN(n29), .Q(next_LO[24]) );
  DFFRX1 \LO_r_reg[23]  ( .D(LO_w[23]), .CK(clk), .RN(n29), .Q(next_LO[23]) );
  DFFRX1 \LO_r_reg[22]  ( .D(LO_w[22]), .CK(clk), .RN(n29), .Q(next_LO[22]) );
  DFFRX1 \LO_r_reg[21]  ( .D(LO_w[21]), .CK(clk), .RN(n29), .Q(next_LO[21]) );
  DFFRX1 \LO_r_reg[20]  ( .D(LO_w[20]), .CK(clk), .RN(n29), .Q(next_LO[20]) );
  DFFRX1 \HI_r_reg[0]  ( .D(HI_w[0]), .CK(clk), .RN(n31), .Q(next_HI[0]) );
  DFFRX1 \LO_r_reg[31]  ( .D(n34), .CK(clk), .RN(n28), .Q(next_LO[31]) );
  DFFRX1 \HI_r_reg[1]  ( .D(HI_w[1]), .CK(clk), .RN(n31), .Q(next_HI[1]) );
  DFFRX1 \HI_r_reg[2]  ( .D(HI_w[2]), .CK(clk), .RN(n31), .Q(next_HI[2]) );
  DFFRX1 \HI_r_reg[3]  ( .D(HI_w[3]), .CK(clk), .RN(n31), .Q(next_HI[3]) );
  DFFRX1 \HI_r_reg[4]  ( .D(HI_w[4]), .CK(clk), .RN(n31), .Q(next_HI[4]) );
  DFFRX1 \HI_r_reg[5]  ( .D(HI_w[5]), .CK(clk), .RN(n31), .Q(next_HI[5]) );
  DFFRX1 \HI_r_reg[6]  ( .D(HI_w[6]), .CK(clk), .RN(n31), .Q(next_HI[6]) );
  DFFRX1 \HI_r_reg[7]  ( .D(HI_w[7]), .CK(clk), .RN(n31), .Q(next_HI[7]) );
  DFFRX1 \HI_r_reg[8]  ( .D(HI_w[8]), .CK(clk), .RN(n31), .Q(next_HI[8]) );
  DFFRX1 \HI_r_reg[9]  ( .D(HI_w[9]), .CK(clk), .RN(n32), .Q(next_HI[9]) );
  DFFRX1 \HI_r_reg[10]  ( .D(HI_w[10]), .CK(clk), .RN(n32), .Q(next_HI[10]) );
  DFFRX1 \HI_r_reg[11]  ( .D(HI_w[11]), .CK(clk), .RN(n32), .Q(next_HI[11]) );
  DFFRX1 \HI_r_reg[12]  ( .D(HI_w[12]), .CK(clk), .RN(n32), .Q(next_HI[12]) );
  DFFRX1 \HI_r_reg[13]  ( .D(HI_w[13]), .CK(clk), .RN(n32), .Q(next_HI[13]) );
  DFFRX1 \HI_r_reg[14]  ( .D(HI_w[14]), .CK(clk), .RN(n32), .Q(next_HI[14]) );
  DFFRX1 \HI_r_reg[15]  ( .D(HI_w[15]), .CK(clk), .RN(n32), .Q(next_HI[15]) );
  DFFRX1 \HI_r_reg[16]  ( .D(HI_w[16]), .CK(clk), .RN(n32), .Q(next_HI[16]) );
  DFFRX1 \HI_r_reg[17]  ( .D(HI_w[17]), .CK(clk), .RN(n32), .Q(next_HI[17]) );
  DFFRX1 \HI_r_reg[18]  ( .D(HI_w[18]), .CK(clk), .RN(n32), .Q(next_HI[18]) );
  DFFRX1 \HI_r_reg[19]  ( .D(HI_w[19]), .CK(clk), .RN(n32), .Q(next_HI[19]) );
  DFFRX1 \HI_r_reg[20]  ( .D(HI_w[20]), .CK(clk), .RN(n32), .Q(next_HI[20]) );
  DFFRX1 \HI_r_reg[21]  ( .D(HI_w[21]), .CK(clk), .RN(n33), .Q(next_HI[21]) );
  DFFRX1 \HI_r_reg[22]  ( .D(HI_w[22]), .CK(clk), .RN(n33), .Q(next_HI[22]) );
  DFFRX1 \HI_r_reg[23]  ( .D(HI_w[23]), .CK(clk), .RN(n33), .Q(next_HI[23]) );
  DFFRX1 \HI_r_reg[24]  ( .D(HI_w[24]), .CK(clk), .RN(n33), .Q(next_HI[24]) );
  DFFRX1 \HI_r_reg[25]  ( .D(HI_w[25]), .CK(clk), .RN(n33), .Q(next_HI[25]) );
  DFFRX1 \HI_r_reg[26]  ( .D(HI_w[26]), .CK(clk), .RN(n33), .Q(next_HI[26]) );
  DFFRX1 \HI_r_reg[27]  ( .D(HI_w[27]), .CK(clk), .RN(n33), .Q(next_HI[27]) );
  DFFRX1 \HI_r_reg[28]  ( .D(HI_w[28]), .CK(clk), .RN(n33), .Q(next_HI[28]) );
  DFFRX1 \HI_r_reg[29]  ( .D(HI_w[29]), .CK(clk), .RN(n33), .Q(next_HI[29]) );
  DFFRX1 \HI_r_reg[30]  ( .D(HI_w[30]), .CK(clk), .RN(n33), .Q(next_HI[30]) );
  DFFRX1 \HI_r_reg[31]  ( .D(HI_w[31]), .CK(clk), .RN(n28), .Q(next_HI[31]) );
  NOR2BX1 U3 ( .AN(n14), .B(n23), .Y(n13) );
  NOR2X1 U4 ( .A(n14), .B(n23), .Y(state_w) );
  CLKBUFX3 U5 ( .A(mul_iter_r[5]), .Y(n23) );
  CLKBUFX3 U8 ( .A(n7), .Y(n5) );
  NOR2X1 U9 ( .A(n5), .B(mul), .Y(n9) );
  CLKBUFX3 U10 ( .A(mul_iter_r[5]), .Y(n24) );
  CLKBUFX3 U11 ( .A(n27), .Y(n32) );
  CLKBUFX3 U12 ( .A(n27), .Y(n31) );
  CLKBUFX3 U13 ( .A(n27), .Y(n30) );
  CLKBUFX3 U14 ( .A(n27), .Y(n29) );
  CLKBUFX3 U15 ( .A(n27), .Y(n28) );
  CLKBUFX3 U16 ( .A(n27), .Y(n33) );
  CLKBUFX3 U17 ( .A(rst), .Y(n27) );
  CLKBUFX3 U18 ( .A(n13), .Y(n3) );
  CLKBUFX3 U19 ( .A(n13), .Y(n4) );
  CLKBUFX3 U20 ( .A(state_w), .Y(n8) );
  CLKBUFX3 U21 ( .A(state_w), .Y(n22) );
  AND2X2 U22 ( .A(multiplicand[1]), .B(next_LO[0]), .Y(N76) );
  AND2X2 U23 ( .A(multiplicand[2]), .B(next_LO[0]), .Y(N77) );
  AND2X2 U24 ( .A(multiplicand[3]), .B(next_LO[0]), .Y(N78) );
  AND2X2 U25 ( .A(multiplicand[4]), .B(next_LO[0]), .Y(N79) );
  AND2X2 U26 ( .A(multiplicand[0]), .B(next_LO[0]), .Y(N75) );
  AO22X1 U27 ( .A0(N74), .A1(n8), .B0(N139), .B1(n3), .Y(HI_w[31]) );
  AO22X1 U28 ( .A0(N73), .A1(n8), .B0(N138), .B1(n3), .Y(HI_w[30]) );
  AO22X1 U29 ( .A0(N72), .A1(n8), .B0(N137), .B1(n3), .Y(HI_w[29]) );
  AO22X1 U30 ( .A0(N71), .A1(n8), .B0(N136), .B1(n3), .Y(HI_w[28]) );
  AO22X1 U31 ( .A0(N70), .A1(n8), .B0(N135), .B1(n3), .Y(HI_w[27]) );
  AND2X2 U32 ( .A(multiplicand[5]), .B(next_LO[0]), .Y(N80) );
  AND2X2 U33 ( .A(multiplicand[6]), .B(next_LO[0]), .Y(N81) );
  AND2X2 U34 ( .A(multiplicand[7]), .B(next_LO[0]), .Y(N82) );
  AND2X2 U35 ( .A(multiplicand[8]), .B(next_LO[0]), .Y(N83) );
  AND2X2 U36 ( .A(multiplicand[9]), .B(next_LO[0]), .Y(N84) );
  AND2X2 U37 ( .A(multiplicand[10]), .B(next_LO[0]), .Y(N85) );
  AND2X2 U38 ( .A(multiplicand[11]), .B(next_LO[0]), .Y(N86) );
  AND2X2 U39 ( .A(multiplicand[12]), .B(next_LO[0]), .Y(N87) );
  AO22X1 U40 ( .A0(N69), .A1(n22), .B0(N134), .B1(n3), .Y(HI_w[26]) );
  AO22X1 U41 ( .A0(N68), .A1(n22), .B0(N133), .B1(n4), .Y(HI_w[25]) );
  AO22X1 U42 ( .A0(N67), .A1(n22), .B0(N132), .B1(n4), .Y(HI_w[24]) );
  AO22X1 U43 ( .A0(N66), .A1(n22), .B0(N131), .B1(n4), .Y(HI_w[23]) );
  AO22X1 U44 ( .A0(N65), .A1(n22), .B0(N130), .B1(n4), .Y(HI_w[22]) );
  AO22X1 U45 ( .A0(N64), .A1(n22), .B0(N129), .B1(n4), .Y(HI_w[21]) );
  AO22X1 U46 ( .A0(N63), .A1(n22), .B0(N128), .B1(n4), .Y(HI_w[20]) );
  AO22X1 U47 ( .A0(N62), .A1(n22), .B0(N127), .B1(n4), .Y(HI_w[19]) );
  AND2X2 U48 ( .A(multiplicand[13]), .B(next_LO[0]), .Y(N88) );
  AND2X2 U49 ( .A(multiplicand[14]), .B(n26), .Y(N89) );
  AND2X2 U50 ( .A(multiplicand[15]), .B(n26), .Y(N90) );
  AND2X2 U51 ( .A(multiplicand[16]), .B(n26), .Y(N91) );
  AND2X2 U52 ( .A(multiplicand[17]), .B(n26), .Y(N92) );
  AND2X2 U53 ( .A(multiplicand[18]), .B(n26), .Y(N93) );
  AND2X2 U54 ( .A(multiplicand[19]), .B(n26), .Y(N94) );
  AND2X2 U55 ( .A(multiplicand[20]), .B(n26), .Y(N95) );
  AO22X1 U56 ( .A0(N54), .A1(n22), .B0(N119), .B1(n4), .Y(HI_w[11]) );
  AO22X1 U57 ( .A0(N61), .A1(n22), .B0(N126), .B1(n4), .Y(HI_w[18]) );
  AO22X1 U58 ( .A0(N60), .A1(n22), .B0(N125), .B1(n4), .Y(HI_w[17]) );
  AO22X1 U59 ( .A0(N59), .A1(n22), .B0(N124), .B1(n4), .Y(HI_w[16]) );
  AO22X1 U60 ( .A0(N58), .A1(n22), .B0(N123), .B1(n4), .Y(HI_w[15]) );
  AO22X1 U61 ( .A0(N57), .A1(n22), .B0(N122), .B1(n4), .Y(HI_w[14]) );
  AO22X1 U62 ( .A0(N56), .A1(n22), .B0(N121), .B1(n4), .Y(HI_w[13]) );
  AO22X1 U63 ( .A0(N55), .A1(n22), .B0(N120), .B1(n4), .Y(HI_w[12]) );
  AND2X2 U64 ( .A(multiplicand[21]), .B(n26), .Y(N96) );
  AND2X2 U65 ( .A(multiplicand[22]), .B(n26), .Y(N97) );
  AND2X2 U66 ( .A(multiplicand[23]), .B(n26), .Y(N98) );
  AND2X2 U67 ( .A(multiplicand[25]), .B(next_LO[0]), .Y(N35) );
  AND2X2 U68 ( .A(multiplicand[26]), .B(next_LO[0]), .Y(N36) );
  AND2X2 U69 ( .A(multiplicand[27]), .B(next_LO[0]), .Y(N37) );
  AND2X2 U70 ( .A(n26), .B(multiplicand[24]), .Y(N99) );
  AO22X1 U71 ( .A0(N53), .A1(n22), .B0(N118), .B1(n4), .Y(HI_w[10]) );
  AO22X1 U72 ( .A0(N52), .A1(n8), .B0(N117), .B1(n3), .Y(HI_w[9]) );
  AO22X1 U73 ( .A0(N51), .A1(n8), .B0(N116), .B1(n3), .Y(HI_w[8]) );
  AO22X1 U74 ( .A0(N50), .A1(n8), .B0(N115), .B1(n3), .Y(HI_w[7]) );
  AO22X1 U75 ( .A0(N49), .A1(n8), .B0(N114), .B1(n3), .Y(HI_w[6]) );
  AO22X1 U76 ( .A0(N48), .A1(n8), .B0(N113), .B1(n3), .Y(HI_w[5]) );
  AO22X1 U77 ( .A0(N47), .A1(n8), .B0(N112), .B1(n3), .Y(HI_w[4]) );
  AND2X2 U78 ( .A(multiplicand[28]), .B(next_LO[0]), .Y(N38) );
  AND2X2 U79 ( .A(multiplicand[29]), .B(next_LO[0]), .Y(N39) );
  AND2X2 U80 ( .A(multiplicand[30]), .B(next_LO[0]), .Y(N40) );
  AND2X2 U81 ( .A(multiplicand[31]), .B(next_LO[0]), .Y(N41) );
  AO22X1 U82 ( .A0(N43), .A1(n22), .B0(N108), .B1(n4), .Y(HI_w[0]) );
  AO22X1 U83 ( .A0(N46), .A1(n8), .B0(N111), .B1(n3), .Y(HI_w[3]) );
  AO22X1 U84 ( .A0(N45), .A1(n8), .B0(N110), .B1(n3), .Y(HI_w[2]) );
  AO22X1 U85 ( .A0(N44), .A1(n22), .B0(N109), .B1(n4), .Y(HI_w[1]) );
  OAI21XL U86 ( .A0(n23), .A1(n11), .B0(n35), .Y(n20) );
  CLKINVX1 U87 ( .A(n9), .Y(n35) );
  NOR2X1 U88 ( .A(N178), .B(n36), .Y(n11) );
  NOR2X1 U89 ( .A(n36), .B(n23), .Y(n10) );
  BUFX4 U90 ( .A(n37), .Y(next_LO[0]) );
  CLKBUFX3 U91 ( .A(n37), .Y(n26) );
  NOR2X1 U92 ( .A(state_r), .B(n36), .Y(mul_stall) );
  CLKINVX1 U93 ( .A(mul), .Y(n36) );
  CLKINVX1 U94 ( .A(n12), .Y(n34) );
  AOI222XL U95 ( .A0(LO[31]), .A1(n23), .B0(N107), .B1(n3), .C0(N42), .C1(n8), 
        .Y(n12) );
  AO22X1 U96 ( .A0(next_LO[2]), .A1(n6), .B0(LO[1]), .B1(n24), .Y(LO_w[1]) );
  AO22X1 U97 ( .A0(next_LO[3]), .A1(n5), .B0(LO[2]), .B1(n23), .Y(LO_w[2]) );
  AO22X1 U98 ( .A0(next_LO[4]), .A1(n5), .B0(LO[3]), .B1(n24), .Y(LO_w[3]) );
  AO22X1 U99 ( .A0(next_LO[5]), .A1(n5), .B0(LO[4]), .B1(n23), .Y(LO_w[4]) );
  AO22X1 U100 ( .A0(next_LO[6]), .A1(n5), .B0(LO[5]), .B1(n23), .Y(LO_w[5]) );
  AO22X1 U101 ( .A0(next_LO[7]), .A1(n5), .B0(LO[6]), .B1(n23), .Y(LO_w[6]) );
  AO22X1 U102 ( .A0(next_LO[8]), .A1(n5), .B0(LO[7]), .B1(n23), .Y(LO_w[7]) );
  AO22X1 U103 ( .A0(next_LO[9]), .A1(n5), .B0(LO[8]), .B1(n23), .Y(LO_w[8]) );
  AO22X1 U104 ( .A0(next_LO[10]), .A1(n5), .B0(LO[9]), .B1(n23), .Y(LO_w[9])
         );
  AO22X1 U105 ( .A0(next_LO[11]), .A1(n6), .B0(LO[10]), .B1(n24), .Y(LO_w[10])
         );
  AO22X1 U106 ( .A0(next_LO[12]), .A1(n6), .B0(LO[11]), .B1(n24), .Y(LO_w[11])
         );
  AO22X1 U107 ( .A0(next_LO[13]), .A1(n6), .B0(LO[12]), .B1(n24), .Y(LO_w[12])
         );
  AO22X1 U108 ( .A0(next_LO[14]), .A1(n6), .B0(LO[13]), .B1(n24), .Y(LO_w[13])
         );
  AO22X1 U109 ( .A0(next_LO[15]), .A1(n6), .B0(LO[14]), .B1(n24), .Y(LO_w[14])
         );
  AO22X1 U110 ( .A0(next_LO[16]), .A1(n6), .B0(LO[15]), .B1(n24), .Y(LO_w[15])
         );
  AO22X1 U111 ( .A0(next_LO[17]), .A1(n6), .B0(LO[16]), .B1(n24), .Y(LO_w[16])
         );
  AO22X1 U112 ( .A0(next_LO[18]), .A1(n6), .B0(LO[17]), .B1(n24), .Y(LO_w[17])
         );
  AO22X1 U113 ( .A0(next_LO[19]), .A1(n6), .B0(LO[18]), .B1(n24), .Y(LO_w[18])
         );
  AO22X1 U114 ( .A0(next_LO[20]), .A1(n6), .B0(LO[19]), .B1(n24), .Y(LO_w[19])
         );
  AO22X1 U115 ( .A0(next_LO[21]), .A1(n5), .B0(LO[20]), .B1(n24), .Y(LO_w[20])
         );
  AO22X1 U116 ( .A0(next_LO[22]), .A1(n5), .B0(LO[21]), .B1(n24), .Y(LO_w[21])
         );
  AO22X1 U117 ( .A0(next_LO[23]), .A1(n5), .B0(LO[22]), .B1(n24), .Y(LO_w[22])
         );
  AO22X1 U118 ( .A0(next_LO[24]), .A1(n5), .B0(LO[23]), .B1(n24), .Y(LO_w[23])
         );
  AO22X1 U119 ( .A0(next_LO[25]), .A1(n5), .B0(LO[24]), .B1(n23), .Y(LO_w[24])
         );
  AO22X1 U120 ( .A0(next_LO[26]), .A1(n5), .B0(LO[25]), .B1(n23), .Y(LO_w[25])
         );
  AO22X1 U121 ( .A0(next_LO[27]), .A1(n5), .B0(LO[26]), .B1(n23), .Y(LO_w[26])
         );
  AO22X1 U122 ( .A0(next_LO[28]), .A1(n5), .B0(LO[27]), .B1(n23), .Y(LO_w[27])
         );
  AO22X1 U123 ( .A0(next_LO[29]), .A1(n5), .B0(LO[28]), .B1(n23), .Y(LO_w[28])
         );
  AO22X1 U124 ( .A0(next_LO[30]), .A1(n5), .B0(LO[29]), .B1(n23), .Y(LO_w[29])
         );
  AO22X1 U125 ( .A0(next_LO[31]), .A1(n5), .B0(LO[30]), .B1(n23), .Y(LO_w[30])
         );
  AO22X1 U126 ( .A0(next_LO[1]), .A1(n6), .B0(LO[0]), .B1(n24), .Y(LO_w[0]) );
  NAND4X1 U127 ( .A(mul_iter_r[4]), .B(mul_iter_r[3]), .C(n15), .D(
        mul_iter_r[2]), .Y(n14) );
  AND2X2 U128 ( .A(mul_iter_r[0]), .B(mul_iter_r[1]), .Y(n15) );
  AO22X1 U129 ( .A0(mul_iter_r[4]), .A1(n9), .B0(N177), .B1(n10), .Y(n19) );
  CLKBUFX3 U130 ( .A(n7), .Y(n6) );
  AO22X1 U131 ( .A0(mul_iter_r[3]), .A1(n9), .B0(N176), .B1(n10), .Y(n18) );
  AO22X1 U132 ( .A0(mul_iter_r[2]), .A1(n9), .B0(N175), .B1(n10), .Y(n17) );
  AO22X1 U133 ( .A0(mul_iter_r[1]), .A1(n9), .B0(N174), .B1(n10), .Y(n16) );
  AO22X1 U134 ( .A0(mul_iter_r[0]), .A1(n9), .B0(N173), .B1(n10), .Y(n21) );
  XOR2X1 U135 ( .A(\add_56/carry[5] ), .B(n24), .Y(N178) );
endmodule


module div_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;
  wire   [32:0] carry;

  ADDFXL U2_30 ( .A(A[30]), .B(n26), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  ADDFXL U2_29 ( .A(A[29]), .B(n24), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  ADDFXL U2_28 ( .A(A[28]), .B(n23), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  ADDFXL U2_27 ( .A(A[27]), .B(n22), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  ADDFXL U2_26 ( .A(A[26]), .B(n21), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  ADDFXL U2_25 ( .A(A[25]), .B(n20), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  ADDFXL U2_24 ( .A(A[24]), .B(n19), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  ADDFXL U2_23 ( .A(A[23]), .B(n18), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  ADDFXL U2_22 ( .A(A[22]), .B(n17), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  ADDFXL U2_21 ( .A(A[21]), .B(n16), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  ADDFXL U2_20 ( .A(A[20]), .B(n15), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  ADDFXL U2_19 ( .A(A[19]), .B(n13), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  ADDFXL U2_18 ( .A(A[18]), .B(n12), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  ADDFXL U2_17 ( .A(A[17]), .B(n11), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  ADDFXL U2_16 ( .A(A[16]), .B(n10), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  ADDFXL U2_15 ( .A(A[15]), .B(n9), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  ADDFXL U2_14 ( .A(A[14]), .B(n8), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFXL U2_13 ( .A(A[13]), .B(n7), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFXL U2_12 ( .A(A[12]), .B(n6), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  ADDFXL U2_11 ( .A(A[11]), .B(n5), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  ADDFXL U2_10 ( .A(A[10]), .B(n4), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  ADDFXL U2_9 ( .A(A[9]), .B(n33), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  ADDFXL U2_8 ( .A(A[8]), .B(n32), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  ADDFXL U2_7 ( .A(A[7]), .B(n31), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  ADDFXL U2_6 ( .A(A[6]), .B(n30), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  ADDFXL U2_5 ( .A(A[5]), .B(n29), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  ADDFXL U2_4 ( .A(A[4]), .B(n28), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFXL U2_3 ( .A(A[3]), .B(n27), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  ADDFXL U2_2 ( .A(A[2]), .B(n25), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  ADDFXL U2_1 ( .A(A[1]), .B(n14), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_31 ( .A(A[31]), .B(n2), .C(carry[31]), .Y(DIFF[31]) );
  CLKINVX1 U1 ( .A(B[0]), .Y(n3) );
  CLKINVX1 U2 ( .A(B[31]), .Y(n2) );
  CLKINVX1 U3 ( .A(B[1]), .Y(n14) );
  NAND2X1 U4 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U5 ( .A(B[2]), .Y(n25) );
  CLKINVX1 U6 ( .A(B[3]), .Y(n27) );
  CLKINVX1 U7 ( .A(B[4]), .Y(n28) );
  CLKINVX1 U8 ( .A(B[5]), .Y(n29) );
  CLKINVX1 U9 ( .A(B[6]), .Y(n30) );
  CLKINVX1 U10 ( .A(B[7]), .Y(n31) );
  CLKINVX1 U11 ( .A(B[8]), .Y(n32) );
  CLKINVX1 U12 ( .A(B[9]), .Y(n33) );
  CLKINVX1 U13 ( .A(B[10]), .Y(n4) );
  CLKINVX1 U14 ( .A(B[11]), .Y(n5) );
  CLKINVX1 U15 ( .A(B[12]), .Y(n6) );
  CLKINVX1 U16 ( .A(B[13]), .Y(n7) );
  CLKINVX1 U17 ( .A(B[14]), .Y(n8) );
  CLKINVX1 U18 ( .A(B[15]), .Y(n9) );
  CLKINVX1 U19 ( .A(B[16]), .Y(n10) );
  CLKINVX1 U20 ( .A(B[17]), .Y(n11) );
  CLKINVX1 U21 ( .A(B[18]), .Y(n12) );
  CLKINVX1 U22 ( .A(B[19]), .Y(n13) );
  CLKINVX1 U23 ( .A(B[20]), .Y(n15) );
  CLKINVX1 U24 ( .A(B[21]), .Y(n16) );
  CLKINVX1 U25 ( .A(B[22]), .Y(n17) );
  CLKINVX1 U26 ( .A(B[23]), .Y(n18) );
  CLKINVX1 U27 ( .A(B[24]), .Y(n19) );
  CLKINVX1 U28 ( .A(B[25]), .Y(n20) );
  CLKINVX1 U29 ( .A(B[26]), .Y(n21) );
  CLKINVX1 U30 ( .A(B[27]), .Y(n22) );
  CLKINVX1 U31 ( .A(B[28]), .Y(n23) );
  CLKINVX1 U32 ( .A(B[29]), .Y(n24) );
  CLKINVX1 U33 ( .A(B[30]), .Y(n26) );
  CLKINVX1 U34 ( .A(A[0]), .Y(n1) );
  XNOR2X1 U35 ( .A(n3), .B(A[0]), .Y(DIFF[0]) );
endmodule


module div_DW01_inc_1 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  ADDHXL U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  ADDHXL U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  ADDHXL U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  ADDHXL U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  ADDHXL U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  ADDHXL U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  ADDHXL U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  ADDHXL U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  ADDHXL U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  ADDHXL U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  ADDHXL U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[31]), .B(A[31]), .Y(SUM[31]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module div_DW01_inc_2 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  ADDHXL U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  ADDHXL U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  ADDHXL U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  ADDHXL U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  ADDHXL U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  ADDHXL U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  ADDHXL U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  ADDHXL U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  ADDHXL U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  ADDHXL U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  ADDHXL U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  ADDHXL U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[31]), .B(A[31]), .Y(SUM[31]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module div_DW01_inc_3 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  ADDHXL U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADDHXL U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  ADDHXL U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  ADDHXL U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  ADDHXL U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  ADDHXL U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  ADDHXL U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  ADDHXL U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  ADDHXL U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  ADDHXL U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  ADDHXL U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[31]), .B(A[31]), .Y(SUM[31]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module div_DW01_inc_4 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  ADDHXL U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADDHXL U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  ADDHXL U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  ADDHXL U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  ADDHXL U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  ADDHXL U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  ADDHXL U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  ADDHXL U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  ADDHXL U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  ADDHXL U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  ADDHXL U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[31]), .B(A[31]), .Y(SUM[31]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module div ( clk, rst, div, divisor, LO, next_HI, next_LO, div_stall );
  input [31:0] divisor;
  input [31:0] LO;
  output [31:0] next_HI;
  output [31:0] next_LO;
  input clk, rst, div;
  output div_stall;
  wire   N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55,
         N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69,
         N70, N71, N72, N73, N108, N109, N110, N111, N112, N113, N114, N115,
         N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N173, N174, N175, N176, N177, N178, N179, N180, N181,
         N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192,
         N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203,
         N204, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258,
         N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269,
         state_r, state_w, N273, N274, N275, N276, N277, N278, n3, n6, n7, n8,
         n9, n11, n12, n13, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n53, n55,
         n57, n59, n61, n63, n65, n68, n70, n72, n74, n76, n78, n80, n82, n84,
         n86, n88, n90, n92, n94, n96, n98, n100, n102, n104, n106, n108, n110,
         n112, n113, n115, n116, n117, n119, n120, n121, n122, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n255,
         n256, n257, n258, n259, n260, \add_130/carry[5] , \add_130/carry[4] ,
         \add_130/carry[3] , \add_130/carry[2] , n2, n4, n5, n10, n14, n36,
         n52, n54, n56, n58, n60, n62, n64, n66, n67, n69, n71, n73, n75, n77,
         n79, n81, n83, n85, n87, n89, n91, n93, n95, n97, n99, n101, n103,
         n105, n107, n109, n111, n114, n118, n123, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287;
  wire   [31:0] HI_r;
  wire   [1:0] sign_r;
  wire   [31:0] divisor_p;
  wire   [5:0] div_iter_r;
  wire   [31:0] diff;
  wire   [31:0] LO_w;
  wire   [31:0] HI_w;

  div_DW01_sub_0 sub_119 ( .A(HI_r), .B(divisor_p), .CI(1'b0), .DIFF(diff) );
  div_DW01_inc_1 add_114 ( .A({n218, n221, n223, n225, n227, n229, n231, n233, 
        n235, n237, n239, n241, n243, n245, n247, n249, n251, n253, n261, n263, 
        n265, n267, n269, n271, n273, n275, n277, n279, n281, n283, n285, n287}), .SUM({N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, 
        N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, 
        N246, N245, N244, N243, N242, N241, N240, N239, N238}) );
  div_DW01_inc_2 add_113 ( .A({n81, n220, n222, n224, n226, n228, n230, n232, 
        n234, n236, n238, n240, n242, n244, n246, n248, n250, n252, n254, n262, 
        n264, n266, n268, n270, n272, n274, n276, n278, n280, n282, n284, n286}), .SUM({N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, 
        N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, 
        N181, N180, N179, N178, N177, N176, N175, N174, N173}) );
  div_DW01_inc_3 add_112 ( .A({n159, n160, n161, n162, n163, n164, n165, n166, 
        n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
        n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190}), .SUM({N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, 
        N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, 
        N116, N115, N114, N113, N112, N111, N110, N109, N108}) );
  div_DW01_inc_4 add_111 ( .A({n127, n128, n129, n130, n131, n132, n133, n134, 
        n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
        n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158}), .SUM({N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45, N44, N43, N42}) );
  DFFRX1 \LO_r_reg[31]  ( .D(LO_w[31]), .CK(clk), .RN(n99), .QN(n159) );
  DFFRX1 \HI_r_reg[31]  ( .D(HI_w[31]), .CK(clk), .RN(n103), .Q(HI_r[31]), 
        .QN(n127) );
  DFFRX1 \LO_r_reg[0]  ( .D(LO_w[0]), .CK(clk), .RN(n93), .QN(n190) );
  ADDHXL \add_130/U1_1_4  ( .A(div_iter_r[4]), .B(\add_130/carry[4] ), .CO(
        \add_130/carry[5] ), .S(N277) );
  ADDHXL \add_130/U1_1_3  ( .A(div_iter_r[3]), .B(\add_130/carry[3] ), .CO(
        \add_130/carry[4] ), .S(N276) );
  ADDHXL \add_130/U1_1_2  ( .A(div_iter_r[2]), .B(\add_130/carry[2] ), .CO(
        \add_130/carry[3] ), .S(N275) );
  ADDHXL \add_130/U1_1_1  ( .A(div_iter_r[1]), .B(div_iter_r[0]), .CO(
        \add_130/carry[2] ), .S(N274) );
  DFFRX1 \HI_r_reg[28]  ( .D(HI_w[28]), .CK(clk), .RN(n103), .Q(HI_r[28]), 
        .QN(n130) );
  DFFRX1 \HI_r_reg[29]  ( .D(HI_w[29]), .CK(clk), .RN(n103), .Q(HI_r[29]), 
        .QN(n129) );
  DFFRX1 \HI_r_reg[30]  ( .D(HI_w[30]), .CK(clk), .RN(n103), .Q(HI_r[30]), 
        .QN(n128) );
  DFFRX1 \LO_r_reg[21]  ( .D(LO_w[21]), .CK(clk), .RN(n97), .QN(n169) );
  DFFRX1 \LO_r_reg[22]  ( .D(LO_w[22]), .CK(clk), .RN(n97), .QN(n168) );
  DFFRX1 \LO_r_reg[23]  ( .D(LO_w[23]), .CK(clk), .RN(n97), .QN(n167) );
  DFFRX1 \LO_r_reg[24]  ( .D(LO_w[24]), .CK(clk), .RN(n97), .QN(n166) );
  DFFRX1 \LO_r_reg[25]  ( .D(LO_w[25]), .CK(clk), .RN(n97), .QN(n165) );
  DFFRX1 \LO_r_reg[26]  ( .D(LO_w[26]), .CK(clk), .RN(n97), .QN(n164) );
  DFFRX1 \LO_r_reg[27]  ( .D(LO_w[27]), .CK(clk), .RN(n97), .QN(n163) );
  DFFRX1 \LO_r_reg[28]  ( .D(LO_w[28]), .CK(clk), .RN(n97), .QN(n162) );
  DFFRX1 \LO_r_reg[29]  ( .D(LO_w[29]), .CK(clk), .RN(n97), .QN(n161) );
  DFFRX1 \LO_r_reg[30]  ( .D(LO_w[30]), .CK(clk), .RN(n99), .QN(n160) );
  DFFRX1 \HI_r_reg[20]  ( .D(HI_w[20]), .CK(clk), .RN(n101), .Q(HI_r[20]), 
        .QN(n138) );
  DFFRX1 \HI_r_reg[21]  ( .D(HI_w[21]), .CK(clk), .RN(n101), .Q(HI_r[21]), 
        .QN(n137) );
  DFFRX1 \HI_r_reg[22]  ( .D(HI_w[22]), .CK(clk), .RN(n103), .Q(HI_r[22]), 
        .QN(n136) );
  DFFRX1 \HI_r_reg[23]  ( .D(HI_w[23]), .CK(clk), .RN(n103), .Q(HI_r[23]), 
        .QN(n135) );
  DFFRX1 \HI_r_reg[24]  ( .D(HI_w[24]), .CK(clk), .RN(n103), .Q(HI_r[24]), 
        .QN(n134) );
  DFFRX1 \HI_r_reg[25]  ( .D(HI_w[25]), .CK(clk), .RN(n103), .Q(HI_r[25]), 
        .QN(n133) );
  DFFRX1 \HI_r_reg[26]  ( .D(HI_w[26]), .CK(clk), .RN(n103), .Q(HI_r[26]), 
        .QN(n132) );
  DFFRX1 \HI_r_reg[27]  ( .D(HI_w[27]), .CK(clk), .RN(n103), .Q(HI_r[27]), 
        .QN(n131) );
  DFFRX1 \LO_r_reg[11]  ( .D(LO_w[11]), .CK(clk), .RN(n95), .QN(n179) );
  DFFRX1 \LO_r_reg[12]  ( .D(LO_w[12]), .CK(clk), .RN(n95), .QN(n178) );
  DFFRX1 \LO_r_reg[13]  ( .D(LO_w[13]), .CK(clk), .RN(n95), .QN(n177) );
  DFFRX1 \LO_r_reg[14]  ( .D(LO_w[14]), .CK(clk), .RN(n95), .QN(n176) );
  DFFRX1 \LO_r_reg[15]  ( .D(LO_w[15]), .CK(clk), .RN(n95), .QN(n175) );
  DFFRX1 \LO_r_reg[16]  ( .D(LO_w[16]), .CK(clk), .RN(n95), .QN(n174) );
  DFFRX1 \LO_r_reg[17]  ( .D(LO_w[17]), .CK(clk), .RN(n95), .QN(n173) );
  DFFRX1 \LO_r_reg[18]  ( .D(LO_w[18]), .CK(clk), .RN(n97), .QN(n172) );
  DFFRX1 \LO_r_reg[19]  ( .D(LO_w[19]), .CK(clk), .RN(n97), .QN(n171) );
  DFFRX1 \LO_r_reg[20]  ( .D(LO_w[20]), .CK(clk), .RN(n97), .QN(n170) );
  DFFRX1 \HI_r_reg[12]  ( .D(HI_w[12]), .CK(clk), .RN(n101), .Q(HI_r[12]), 
        .QN(n146) );
  DFFRX1 \HI_r_reg[13]  ( .D(HI_w[13]), .CK(clk), .RN(n101), .Q(HI_r[13]), 
        .QN(n145) );
  DFFRX1 \HI_r_reg[14]  ( .D(HI_w[14]), .CK(clk), .RN(n101), .Q(HI_r[14]), 
        .QN(n144) );
  DFFRX1 \HI_r_reg[15]  ( .D(HI_w[15]), .CK(clk), .RN(n101), .Q(HI_r[15]), 
        .QN(n143) );
  DFFRX1 \HI_r_reg[16]  ( .D(HI_w[16]), .CK(clk), .RN(n101), .Q(HI_r[16]), 
        .QN(n142) );
  DFFRX1 \HI_r_reg[17]  ( .D(HI_w[17]), .CK(clk), .RN(n101), .Q(HI_r[17]), 
        .QN(n141) );
  DFFRX1 \HI_r_reg[18]  ( .D(HI_w[18]), .CK(clk), .RN(n101), .Q(HI_r[18]), 
        .QN(n140) );
  DFFRX1 \HI_r_reg[19]  ( .D(HI_w[19]), .CK(clk), .RN(n101), .Q(HI_r[19]), 
        .QN(n139) );
  DFFRX1 \LO_r_reg[2]  ( .D(LO_w[2]), .CK(clk), .RN(n93), .QN(n188) );
  DFFRX1 \LO_r_reg[3]  ( .D(LO_w[3]), .CK(clk), .RN(n93), .QN(n187) );
  DFFRX1 \LO_r_reg[4]  ( .D(LO_w[4]), .CK(clk), .RN(n93), .QN(n186) );
  DFFRX1 \LO_r_reg[5]  ( .D(LO_w[5]), .CK(clk), .RN(n93), .QN(n185) );
  DFFRX1 \LO_r_reg[6]  ( .D(LO_w[6]), .CK(clk), .RN(n95), .QN(n184) );
  DFFRX1 \LO_r_reg[7]  ( .D(LO_w[7]), .CK(clk), .RN(n95), .QN(n183) );
  DFFRX1 \LO_r_reg[8]  ( .D(LO_w[8]), .CK(clk), .RN(n95), .QN(n182) );
  DFFRX1 \LO_r_reg[9]  ( .D(LO_w[9]), .CK(clk), .RN(n95), .QN(n181) );
  DFFRX1 \LO_r_reg[10]  ( .D(LO_w[10]), .CK(clk), .RN(n95), .QN(n180) );
  DFFRX1 \HI_r_reg[4]  ( .D(HI_w[4]), .CK(clk), .RN(n99), .Q(HI_r[4]), .QN(
        n154) );
  DFFRX1 \HI_r_reg[5]  ( .D(HI_w[5]), .CK(clk), .RN(n99), .Q(HI_r[5]), .QN(
        n153) );
  DFFRX1 \HI_r_reg[6]  ( .D(HI_w[6]), .CK(clk), .RN(n99), .Q(HI_r[6]), .QN(
        n152) );
  DFFRX1 \HI_r_reg[7]  ( .D(HI_w[7]), .CK(clk), .RN(n99), .Q(HI_r[7]), .QN(
        n151) );
  DFFRX1 \HI_r_reg[8]  ( .D(HI_w[8]), .CK(clk), .RN(n99), .Q(HI_r[8]), .QN(
        n150) );
  DFFRX1 \HI_r_reg[9]  ( .D(HI_w[9]), .CK(clk), .RN(n99), .Q(HI_r[9]), .QN(
        n149) );
  DFFRX1 \HI_r_reg[10]  ( .D(HI_w[10]), .CK(clk), .RN(n101), .Q(HI_r[10]), 
        .QN(n148) );
  DFFRX1 \HI_r_reg[11]  ( .D(HI_w[11]), .CK(clk), .RN(n101), .Q(HI_r[11]), 
        .QN(n147) );
  DFFRX1 \HI_r_reg[1]  ( .D(HI_w[1]), .CK(clk), .RN(n99), .Q(HI_r[1]), .QN(
        n157) );
  DFFRX1 \HI_r_reg[2]  ( .D(HI_w[2]), .CK(clk), .RN(n99), .Q(HI_r[2]), .QN(
        n156) );
  DFFRX1 \HI_r_reg[3]  ( .D(HI_w[3]), .CK(clk), .RN(n99), .Q(HI_r[3]), .QN(
        n155) );
  DFFRX1 \HI_r_reg[0]  ( .D(HI_w[0]), .CK(clk), .RN(n99), .Q(HI_r[0]), .QN(
        n158) );
  DFFRX1 \LO_r_reg[1]  ( .D(LO_w[1]), .CK(clk), .RN(n93), .QN(n189) );
  DFFRX1 state_r_reg ( .D(state_w), .CK(clk), .RN(n93), .Q(state_r) );
  DFFRX1 \sign_r_reg[0]  ( .D(n124), .CK(clk), .RN(n103), .Q(sign_r[0]) );
  DFFRX1 \sign_r_reg[1]  ( .D(n125), .CK(clk), .RN(n103), .Q(sign_r[1]) );
  DFFRX1 \div_iter_r_reg[3]  ( .D(n257), .CK(clk), .RN(n93), .Q(div_iter_r[3]), 
        .QN(n120) );
  DFFRX1 \div_iter_r_reg[2]  ( .D(n256), .CK(clk), .RN(n93), .Q(div_iter_r[2]), 
        .QN(n121) );
  DFFRX1 \div_iter_r_reg[1]  ( .D(n255), .CK(clk), .RN(n93), .Q(div_iter_r[1]), 
        .QN(n122) );
  DFFRX1 \div_iter_r_reg[0]  ( .D(n260), .CK(clk), .RN(n93), .Q(div_iter_r[0]), 
        .QN(N273) );
  DFFRX1 \div_iter_r_reg[4]  ( .D(n258), .CK(clk), .RN(n93), .Q(div_iter_r[4]), 
        .QN(n119) );
  DFFSX2 \div_iter_r_reg[5]  ( .D(n259), .CK(clk), .SN(rst), .Q(div_iter_r[5]), 
        .QN(n126) );
  NAND2X1 U3 ( .A(state_w), .B(n107), .Y(n51) );
  NAND2X1 U4 ( .A(n113), .B(n107), .Y(n39) );
  CLKINVX1 U5 ( .A(n113), .Y(n217) );
  NAND2X1 U6 ( .A(n113), .B(diff[31]), .Y(n34) );
  NAND2X1 U7 ( .A(diff[31]), .B(state_w), .Y(n40) );
  NAND2X1 U8 ( .A(div_iter_r[5]), .B(n218), .Y(n12) );
  NOR2X1 U9 ( .A(n218), .B(n126), .Y(n6) );
  XOR2X1 U11 ( .A(sign_r[0]), .B(n77), .Y(n3) );
  CLKBUFX3 U12 ( .A(sign_r[1]), .Y(n79) );
  CLKBUFX3 U13 ( .A(sign_r[1]), .Y(n75) );
  CLKBUFX3 U14 ( .A(n89), .Y(n103) );
  CLKBUFX3 U15 ( .A(n89), .Y(n101) );
  CLKBUFX3 U16 ( .A(n91), .Y(n99) );
  CLKBUFX3 U17 ( .A(n91), .Y(n97) );
  CLKBUFX3 U18 ( .A(n89), .Y(n95) );
  CLKBUFX3 U19 ( .A(n91), .Y(n93) );
  CLKBUFX3 U20 ( .A(rst), .Y(n89) );
  CLKBUFX3 U21 ( .A(rst), .Y(n91) );
  INVX3 U22 ( .A(divisor[31]), .Y(n81) );
  CLKBUFX3 U23 ( .A(n11), .Y(n64) );
  INVX3 U24 ( .A(divisor[31]), .Y(n83) );
  AND2X2 U25 ( .A(n10), .B(n40), .Y(n11) );
  CLKBUFX3 U26 ( .A(n51), .Y(n5) );
  CLKBUFX3 U27 ( .A(divisor[31]), .Y(n85) );
  CLKBUFX3 U28 ( .A(divisor[31]), .Y(n87) );
  CLKBUFX3 U29 ( .A(n39), .Y(n52) );
  CLKBUFX3 U30 ( .A(n39), .Y(n54) );
  CLKBUFX3 U31 ( .A(n51), .Y(n10) );
  CLKBUFX3 U32 ( .A(n217), .Y(n2) );
  CLKBUFX3 U33 ( .A(n217), .Y(n4) );
  CLKBUFX3 U34 ( .A(n40), .Y(n14) );
  CLKBUFX3 U35 ( .A(n40), .Y(n36) );
  CLKBUFX3 U36 ( .A(n34), .Y(n56) );
  CLKBUFX3 U37 ( .A(n34), .Y(n58) );
  CLKBUFX3 U38 ( .A(n12), .Y(n60) );
  CLKBUFX3 U39 ( .A(n12), .Y(n62) );
  CLKBUFX3 U40 ( .A(n3), .Y(n69) );
  CLKBUFX3 U41 ( .A(n3), .Y(n71) );
  CLKBUFX3 U42 ( .A(n3), .Y(n73) );
  OAI211X1 U43 ( .A0(n190), .A1(n56), .B0(n35), .C0(n105), .Y(LO_w[1]) );
  NAND2X1 U44 ( .A(N238), .B(n67), .Y(n35) );
  CLKINVX1 U45 ( .A(n37), .Y(n105) );
  CLKINVX1 U46 ( .A(divisor[0]), .Y(n286) );
  CLKINVX1 U47 ( .A(divisor[1]), .Y(n284) );
  CLKINVX1 U48 ( .A(divisor[2]), .Y(n282) );
  CLKINVX1 U49 ( .A(divisor[3]), .Y(n280) );
  CLKINVX1 U50 ( .A(divisor[4]), .Y(n278) );
  CLKINVX1 U51 ( .A(divisor[5]), .Y(n276) );
  CLKINVX1 U52 ( .A(divisor[6]), .Y(n274) );
  CLKINVX1 U53 ( .A(divisor[7]), .Y(n272) );
  OAI21XL U54 ( .A0(n190), .A1(n14), .B0(n5), .Y(LO_w[0]) );
  CLKINVX1 U55 ( .A(diff[31]), .Y(n107) );
  AO22X1 U56 ( .A0(n81), .A1(divisor[0]), .B0(N173), .B1(n87), .Y(divisor_p[0]) );
  CLKINVX1 U57 ( .A(divisor[8]), .Y(n270) );
  CLKINVX1 U58 ( .A(divisor[9]), .Y(n268) );
  CLKINVX1 U59 ( .A(divisor[10]), .Y(n266) );
  CLKINVX1 U60 ( .A(divisor[11]), .Y(n264) );
  CLKINVX1 U61 ( .A(divisor[12]), .Y(n262) );
  CLKINVX1 U62 ( .A(divisor[13]), .Y(n254) );
  CLKINVX1 U63 ( .A(divisor[14]), .Y(n252) );
  CLKINVX1 U64 ( .A(divisor[15]), .Y(n250) );
  CLKINVX1 U65 ( .A(divisor[16]), .Y(n248) );
  CLKINVX1 U66 ( .A(divisor[17]), .Y(n246) );
  CLKINVX1 U67 ( .A(divisor[18]), .Y(n244) );
  CLKINVX1 U68 ( .A(divisor[19]), .Y(n242) );
  CLKINVX1 U69 ( .A(divisor[20]), .Y(n240) );
  CLKINVX1 U70 ( .A(divisor[21]), .Y(n238) );
  CLKINVX1 U71 ( .A(divisor[22]), .Y(n236) );
  CLKINVX1 U72 ( .A(divisor[23]), .Y(n234) );
  CLKINVX1 U73 ( .A(divisor[24]), .Y(n232) );
  CLKINVX1 U74 ( .A(divisor[25]), .Y(n230) );
  CLKINVX1 U75 ( .A(divisor[26]), .Y(n228) );
  CLKINVX1 U76 ( .A(divisor[27]), .Y(n226) );
  CLKINVX1 U77 ( .A(divisor[28]), .Y(n224) );
  CLKINVX1 U78 ( .A(divisor[29]), .Y(n222) );
  CLKINVX1 U79 ( .A(divisor[30]), .Y(n220) );
  CLKINVX1 U80 ( .A(diff[30]), .Y(n109) );
  CLKINVX1 U81 ( .A(diff[29]), .Y(n111) );
  CLKINVX1 U82 ( .A(diff[28]), .Y(n114) );
  CLKINVX1 U83 ( .A(diff[27]), .Y(n118) );
  CLKINVX1 U84 ( .A(diff[26]), .Y(n123) );
  CLKINVX1 U85 ( .A(diff[25]), .Y(n191) );
  CLKINVX1 U86 ( .A(LO[0]), .Y(n287) );
  CLKINVX1 U87 ( .A(LO[1]), .Y(n285) );
  CLKINVX1 U88 ( .A(LO[24]), .Y(n233) );
  CLKINVX1 U89 ( .A(LO[2]), .Y(n283) );
  CLKINVX1 U90 ( .A(LO[3]), .Y(n281) );
  CLKINVX1 U91 ( .A(LO[4]), .Y(n279) );
  CLKINVX1 U92 ( .A(LO[5]), .Y(n277) );
  CLKINVX1 U93 ( .A(LO[6]), .Y(n275) );
  CLKINVX1 U94 ( .A(LO[7]), .Y(n273) );
  CLKINVX1 U95 ( .A(LO[8]), .Y(n271) );
  CLKINVX1 U96 ( .A(LO[9]), .Y(n269) );
  CLKINVX1 U97 ( .A(LO[10]), .Y(n267) );
  CLKINVX1 U98 ( .A(LO[11]), .Y(n265) );
  CLKINVX1 U99 ( .A(LO[12]), .Y(n263) );
  CLKINVX1 U100 ( .A(LO[13]), .Y(n261) );
  CLKINVX1 U101 ( .A(LO[14]), .Y(n253) );
  CLKINVX1 U102 ( .A(LO[15]), .Y(n251) );
  CLKINVX1 U103 ( .A(LO[16]), .Y(n249) );
  CLKINVX1 U104 ( .A(LO[17]), .Y(n247) );
  CLKINVX1 U105 ( .A(LO[18]), .Y(n245) );
  CLKINVX1 U106 ( .A(LO[19]), .Y(n243) );
  CLKINVX1 U107 ( .A(LO[20]), .Y(n241) );
  CLKINVX1 U108 ( .A(LO[21]), .Y(n239) );
  CLKINVX1 U109 ( .A(LO[22]), .Y(n237) );
  CLKINVX1 U110 ( .A(LO[23]), .Y(n235) );
  CLKINVX1 U111 ( .A(LO[25]), .Y(n231) );
  CLKINVX1 U112 ( .A(LO[26]), .Y(n229) );
  CLKINVX1 U113 ( .A(LO[27]), .Y(n227) );
  CLKINVX1 U114 ( .A(LO[28]), .Y(n225) );
  CLKINVX1 U115 ( .A(LO[29]), .Y(n223) );
  CLKINVX1 U116 ( .A(diff[24]), .Y(n192) );
  CLKINVX1 U117 ( .A(diff[23]), .Y(n193) );
  CLKINVX1 U118 ( .A(diff[22]), .Y(n194) );
  CLKINVX1 U119 ( .A(diff[21]), .Y(n195) );
  CLKINVX1 U120 ( .A(diff[20]), .Y(n196) );
  CLKINVX1 U121 ( .A(diff[19]), .Y(n197) );
  CLKINVX1 U122 ( .A(diff[18]), .Y(n198) );
  CLKINVX1 U123 ( .A(diff[17]), .Y(n199) );
  CLKINVX1 U124 ( .A(LO[30]), .Y(n221) );
  CLKINVX1 U125 ( .A(diff[16]), .Y(n200) );
  CLKINVX1 U126 ( .A(diff[15]), .Y(n201) );
  CLKINVX1 U127 ( .A(diff[14]), .Y(n202) );
  CLKINVX1 U128 ( .A(diff[13]), .Y(n203) );
  CLKINVX1 U129 ( .A(diff[12]), .Y(n204) );
  CLKINVX1 U130 ( .A(diff[11]), .Y(n205) );
  CLKINVX1 U131 ( .A(diff[10]), .Y(n206) );
  CLKINVX1 U132 ( .A(diff[9]), .Y(n207) );
  CLKINVX1 U133 ( .A(diff[7]), .Y(n209) );
  CLKINVX1 U134 ( .A(diff[6]), .Y(n210) );
  CLKINVX1 U135 ( .A(diff[5]), .Y(n211) );
  CLKINVX1 U136 ( .A(diff[4]), .Y(n212) );
  CLKINVX1 U137 ( .A(diff[3]), .Y(n213) );
  CLKINVX1 U138 ( .A(diff[2]), .Y(n214) );
  CLKINVX1 U139 ( .A(diff[1]), .Y(n215) );
  CLKINVX1 U140 ( .A(diff[8]), .Y(n208) );
  CLKINVX1 U141 ( .A(LO[31]), .Y(n218) );
  CLKBUFX3 U142 ( .A(n6), .Y(n66) );
  CLKBUFX3 U143 ( .A(n6), .Y(n67) );
  NOR2BX1 U144 ( .AN(n116), .B(div_iter_r[5]), .Y(state_w) );
  NOR2X1 U145 ( .A(div_iter_r[5]), .B(n116), .Y(n113) );
  NAND2X1 U146 ( .A(n219), .B(div_iter_r[5]), .Y(n7) );
  NOR2X1 U147 ( .A(n219), .B(div_iter_r[5]), .Y(n8) );
  OAI222XL U148 ( .A0(n128), .A1(n56), .B0(n52), .B1(n109), .C0(n127), .C1(n14), .Y(HI_w[31]) );
  OAI221XL U149 ( .A0(n62), .A1(n287), .B0(n38), .B1(n189), .C0(n52), .Y(n37)
         );
  OA21XL U150 ( .A0(diff[31]), .A1(div_iter_r[5]), .B0(n40), .Y(n38) );
  OAI221XL U151 ( .A0(n128), .A1(n36), .B0(n5), .B1(n109), .C0(n68), .Y(
        HI_w[30]) );
  OA22X1 U152 ( .A0(n58), .A1(n129), .B0(n111), .B1(n54), .Y(n68) );
  OAI221XL U153 ( .A0(n129), .A1(n36), .B0(n5), .B1(n111), .C0(n72), .Y(
        HI_w[29]) );
  OA22X1 U154 ( .A0(n58), .A1(n130), .B0(n114), .B1(n54), .Y(n72) );
  OAI221XL U155 ( .A0(n130), .A1(n36), .B0(n5), .B1(n114), .C0(n74), .Y(
        HI_w[28]) );
  OA22X1 U156 ( .A0(n58), .A1(n131), .B0(n118), .B1(n54), .Y(n74) );
  OAI221XL U157 ( .A0(n131), .A1(n36), .B0(n5), .B1(n118), .C0(n76), .Y(
        HI_w[27]) );
  OA22X1 U158 ( .A0(n58), .A1(n132), .B0(n123), .B1(n54), .Y(n76) );
  OAI221XL U159 ( .A0(n132), .A1(n36), .B0(n5), .B1(n123), .C0(n78), .Y(
        HI_w[26]) );
  OA22X1 U160 ( .A0(n58), .A1(n133), .B0(n191), .B1(n54), .Y(n78) );
  OAI221XL U161 ( .A0(n133), .A1(n36), .B0(n5), .B1(n191), .C0(n80), .Y(
        HI_w[25]) );
  OA22X1 U162 ( .A0(n58), .A1(n134), .B0(n192), .B1(n54), .Y(n80) );
  OAI221XL U163 ( .A0(n134), .A1(n36), .B0(n10), .B1(n192), .C0(n82), .Y(
        HI_w[24]) );
  OA22X1 U164 ( .A0(n58), .A1(n135), .B0(n193), .B1(n54), .Y(n82) );
  OAI221XL U165 ( .A0(n135), .A1(n36), .B0(n51), .B1(n193), .C0(n84), .Y(
        HI_w[23]) );
  OA22X1 U166 ( .A0(n58), .A1(n136), .B0(n194), .B1(n54), .Y(n84) );
  OAI221XL U167 ( .A0(n136), .A1(n14), .B0(n51), .B1(n194), .C0(n86), .Y(
        HI_w[22]) );
  OA22X1 U168 ( .A0(n58), .A1(n137), .B0(n195), .B1(n54), .Y(n86) );
  OAI221XL U169 ( .A0(n137), .A1(n14), .B0(n5), .B1(n195), .C0(n88), .Y(
        HI_w[21]) );
  OA22X1 U170 ( .A0(n58), .A1(n138), .B0(n196), .B1(n52), .Y(n88) );
  OAI221XL U171 ( .A0(n138), .A1(n14), .B0(n5), .B1(n196), .C0(n90), .Y(
        HI_w[20]) );
  OA22X1 U172 ( .A0(n56), .A1(n139), .B0(n197), .B1(n52), .Y(n90) );
  OAI221XL U173 ( .A0(n139), .A1(n14), .B0(n5), .B1(n197), .C0(n94), .Y(
        HI_w[19]) );
  OA22X1 U174 ( .A0(n56), .A1(n140), .B0(n198), .B1(n52), .Y(n94) );
  OAI221XL U175 ( .A0(n140), .A1(n14), .B0(n5), .B1(n198), .C0(n96), .Y(
        HI_w[18]) );
  OA22X1 U176 ( .A0(n56), .A1(n141), .B0(n199), .B1(n52), .Y(n96) );
  OAI221XL U177 ( .A0(n141), .A1(n14), .B0(n5), .B1(n199), .C0(n98), .Y(
        HI_w[17]) );
  OA22X1 U178 ( .A0(n56), .A1(n142), .B0(n200), .B1(n52), .Y(n98) );
  OAI221XL U179 ( .A0(n142), .A1(n14), .B0(n5), .B1(n200), .C0(n100), .Y(
        HI_w[16]) );
  OA22X1 U180 ( .A0(n56), .A1(n143), .B0(n201), .B1(n52), .Y(n100) );
  OAI221XL U181 ( .A0(n143), .A1(n14), .B0(n5), .B1(n201), .C0(n102), .Y(
        HI_w[15]) );
  OA22X1 U182 ( .A0(n56), .A1(n144), .B0(n202), .B1(n52), .Y(n102) );
  OAI221XL U183 ( .A0(n144), .A1(n14), .B0(n5), .B1(n202), .C0(n104), .Y(
        HI_w[14]) );
  OA22X1 U184 ( .A0(n56), .A1(n145), .B0(n203), .B1(n52), .Y(n104) );
  OAI221XL U185 ( .A0(n145), .A1(n14), .B0(n5), .B1(n203), .C0(n106), .Y(
        HI_w[13]) );
  OA22X1 U186 ( .A0(n56), .A1(n146), .B0(n204), .B1(n52), .Y(n106) );
  OAI221XL U187 ( .A0(n146), .A1(n14), .B0(n5), .B1(n204), .C0(n108), .Y(
        HI_w[12]) );
  OA22X1 U188 ( .A0(n56), .A1(n147), .B0(n205), .B1(n52), .Y(n108) );
  OAI221XL U189 ( .A0(n147), .A1(n14), .B0(n5), .B1(n205), .C0(n110), .Y(
        HI_w[11]) );
  OA22X1 U190 ( .A0(n56), .A1(n148), .B0(n206), .B1(n52), .Y(n110) );
  OAI221XL U191 ( .A0(n148), .A1(n14), .B0(n5), .B1(n206), .C0(n112), .Y(
        HI_w[10]) );
  OA22X1 U192 ( .A0(n58), .A1(n149), .B0(n207), .B1(n54), .Y(n112) );
  OAI221XL U193 ( .A0(n152), .A1(n36), .B0(n10), .B1(n210), .C0(n59), .Y(
        HI_w[6]) );
  OA22X1 U194 ( .A0(n56), .A1(n153), .B0(n211), .B1(n54), .Y(n59) );
  OAI221XL U195 ( .A0(n153), .A1(n36), .B0(n51), .B1(n211), .C0(n61), .Y(
        HI_w[5]) );
  OA22X1 U196 ( .A0(n58), .A1(n154), .B0(n212), .B1(n54), .Y(n61) );
  OAI221XL U197 ( .A0(n154), .A1(n36), .B0(n51), .B1(n212), .C0(n63), .Y(
        HI_w[4]) );
  OA22X1 U198 ( .A0(n58), .A1(n155), .B0(n213), .B1(n54), .Y(n63) );
  OAI221XL U199 ( .A0(n155), .A1(n36), .B0(n10), .B1(n213), .C0(n65), .Y(
        HI_w[3]) );
  OA22X1 U200 ( .A0(n58), .A1(n156), .B0(n214), .B1(n54), .Y(n65) );
  OAI221XL U201 ( .A0(n156), .A1(n36), .B0(n10), .B1(n214), .C0(n70), .Y(
        HI_w[2]) );
  OA22X1 U202 ( .A0(n58), .A1(n157), .B0(n215), .B1(n54), .Y(n70) );
  OAI221XL U203 ( .A0(n157), .A1(n14), .B0(n5), .B1(n215), .C0(n92), .Y(
        HI_w[1]) );
  OA22X1 U204 ( .A0(n56), .A1(n158), .B0(n216), .B1(n52), .Y(n92) );
  OAI221XL U205 ( .A0(n158), .A1(n36), .B0(n10), .B1(n216), .C0(n115), .Y(
        HI_w[0]) );
  AOI2BB2X1 U206 ( .B0(N269), .B1(n67), .A0N(n159), .A1N(n2), .Y(n115) );
  OAI221XL U207 ( .A0(n159), .A1(n64), .B0(n221), .B1(n60), .C0(n21), .Y(
        LO_w[31]) );
  AOI2BB2X1 U208 ( .B0(N268), .B1(n67), .A0N(n160), .A1N(n4), .Y(n21) );
  OAI221XL U209 ( .A0(n160), .A1(n11), .B0(n223), .B1(n60), .C0(n22), .Y(
        LO_w[30]) );
  AOI2BB2X1 U210 ( .B0(N267), .B1(n67), .A0N(n161), .A1N(n4), .Y(n22) );
  OAI221XL U211 ( .A0(n161), .A1(n11), .B0(n225), .B1(n60), .C0(n24), .Y(
        LO_w[29]) );
  AOI2BB2X1 U212 ( .B0(N266), .B1(n67), .A0N(n162), .A1N(n4), .Y(n24) );
  OAI221XL U213 ( .A0(n162), .A1(n11), .B0(n227), .B1(n60), .C0(n25), .Y(
        LO_w[28]) );
  AOI2BB2X1 U214 ( .B0(N265), .B1(n66), .A0N(n163), .A1N(n4), .Y(n25) );
  OAI221XL U215 ( .A0(n163), .A1(n11), .B0(n229), .B1(n60), .C0(n26), .Y(
        LO_w[27]) );
  AOI2BB2X1 U216 ( .B0(N264), .B1(n67), .A0N(n164), .A1N(n4), .Y(n26) );
  OAI221XL U217 ( .A0(n164), .A1(n11), .B0(n231), .B1(n60), .C0(n27), .Y(
        LO_w[26]) );
  AOI2BB2X1 U218 ( .B0(N263), .B1(n66), .A0N(n165), .A1N(n4), .Y(n27) );
  OAI221XL U219 ( .A0(n165), .A1(n11), .B0(n233), .B1(n62), .C0(n28), .Y(
        LO_w[25]) );
  AOI2BB2X1 U220 ( .B0(N262), .B1(n67), .A0N(n166), .A1N(n4), .Y(n28) );
  OAI221XL U221 ( .A0(n166), .A1(n11), .B0(n235), .B1(n60), .C0(n29), .Y(
        LO_w[24]) );
  AOI2BB2X1 U222 ( .B0(N261), .B1(n66), .A0N(n167), .A1N(n4), .Y(n29) );
  OAI221XL U223 ( .A0(n167), .A1(n11), .B0(n237), .B1(n12), .C0(n30), .Y(
        LO_w[23]) );
  AOI2BB2X1 U224 ( .B0(N260), .B1(n67), .A0N(n168), .A1N(n4), .Y(n30) );
  OAI221XL U225 ( .A0(n168), .A1(n64), .B0(n239), .B1(n12), .C0(n31), .Y(
        LO_w[22]) );
  AOI2BB2X1 U226 ( .B0(N259), .B1(n66), .A0N(n169), .A1N(n4), .Y(n31) );
  OAI221XL U227 ( .A0(n169), .A1(n64), .B0(n241), .B1(n60), .C0(n32), .Y(
        LO_w[21]) );
  AOI2BB2X1 U228 ( .B0(N258), .B1(n66), .A0N(n170), .A1N(n2), .Y(n32) );
  OAI221XL U229 ( .A0(n170), .A1(n64), .B0(n243), .B1(n60), .C0(n33), .Y(
        LO_w[20]) );
  AOI2BB2X1 U230 ( .B0(N257), .B1(n66), .A0N(n171), .A1N(n2), .Y(n33) );
  OAI221XL U231 ( .A0(n171), .A1(n64), .B0(n245), .B1(n60), .C0(n41), .Y(
        LO_w[19]) );
  AOI2BB2X1 U232 ( .B0(N256), .B1(n66), .A0N(n172), .A1N(n2), .Y(n41) );
  OAI221XL U233 ( .A0(n172), .A1(n64), .B0(n247), .B1(n60), .C0(n42), .Y(
        LO_w[18]) );
  AOI2BB2X1 U234 ( .B0(N255), .B1(n66), .A0N(n173), .A1N(n2), .Y(n42) );
  OAI221XL U235 ( .A0(n173), .A1(n64), .B0(n249), .B1(n60), .C0(n43), .Y(
        LO_w[17]) );
  AOI2BB2X1 U236 ( .B0(N254), .B1(n66), .A0N(n174), .A1N(n2), .Y(n43) );
  OAI221XL U237 ( .A0(n174), .A1(n64), .B0(n251), .B1(n60), .C0(n44), .Y(
        LO_w[16]) );
  AOI2BB2X1 U238 ( .B0(N253), .B1(n66), .A0N(n175), .A1N(n2), .Y(n44) );
  OAI221XL U239 ( .A0(n175), .A1(n64), .B0(n253), .B1(n60), .C0(n45), .Y(
        LO_w[15]) );
  AOI2BB2X1 U240 ( .B0(N252), .B1(n66), .A0N(n176), .A1N(n2), .Y(n45) );
  OAI221XL U241 ( .A0(n176), .A1(n64), .B0(n261), .B1(n60), .C0(n46), .Y(
        LO_w[14]) );
  AOI2BB2X1 U242 ( .B0(N251), .B1(n66), .A0N(n177), .A1N(n2), .Y(n46) );
  OAI221XL U243 ( .A0(n177), .A1(n64), .B0(n263), .B1(n60), .C0(n47), .Y(
        LO_w[13]) );
  AOI2BB2X1 U244 ( .B0(N250), .B1(n66), .A0N(n178), .A1N(n2), .Y(n47) );
  OAI221XL U245 ( .A0(n178), .A1(n64), .B0(n265), .B1(n60), .C0(n48), .Y(
        LO_w[12]) );
  AOI2BB2X1 U246 ( .B0(N249), .B1(n66), .A0N(n179), .A1N(n2), .Y(n48) );
  OAI221XL U247 ( .A0(n179), .A1(n64), .B0(n267), .B1(n60), .C0(n49), .Y(
        LO_w[11]) );
  AOI2BB2X1 U248 ( .B0(N248), .B1(n66), .A0N(n180), .A1N(n2), .Y(n49) );
  OAI221XL U249 ( .A0(n180), .A1(n64), .B0(n269), .B1(n12), .C0(n50), .Y(
        LO_w[10]) );
  AOI2BB2X1 U250 ( .B0(N247), .B1(n66), .A0N(n181), .A1N(n2), .Y(n50) );
  OAI221XL U251 ( .A0(n181), .A1(n64), .B0(n271), .B1(n60), .C0(n13), .Y(
        LO_w[9]) );
  AOI2BB2X1 U252 ( .B0(N246), .B1(n67), .A0N(n182), .A1N(n2), .Y(n13) );
  OAI221XL U253 ( .A0(n182), .A1(n11), .B0(n273), .B1(n62), .C0(n15), .Y(
        LO_w[8]) );
  AOI2BB2X1 U254 ( .B0(N245), .B1(n67), .A0N(n183), .A1N(n4), .Y(n15) );
  OAI221XL U255 ( .A0(n183), .A1(n11), .B0(n275), .B1(n62), .C0(n16), .Y(
        LO_w[7]) );
  AOI2BB2X1 U256 ( .B0(N244), .B1(n67), .A0N(n184), .A1N(n2), .Y(n16) );
  OAI221XL U257 ( .A0(n184), .A1(n11), .B0(n277), .B1(n62), .C0(n17), .Y(
        LO_w[6]) );
  AOI2BB2X1 U258 ( .B0(N243), .B1(n67), .A0N(n185), .A1N(n4), .Y(n17) );
  OAI221XL U259 ( .A0(n185), .A1(n11), .B0(n279), .B1(n62), .C0(n18), .Y(
        LO_w[5]) );
  AOI2BB2X1 U260 ( .B0(N242), .B1(n67), .A0N(n186), .A1N(n217), .Y(n18) );
  OAI221XL U261 ( .A0(n186), .A1(n64), .B0(n281), .B1(n62), .C0(n19), .Y(
        LO_w[4]) );
  AOI2BB2X1 U262 ( .B0(N241), .B1(n67), .A0N(n187), .A1N(n4), .Y(n19) );
  OAI221XL U263 ( .A0(n187), .A1(n64), .B0(n283), .B1(n62), .C0(n20), .Y(
        LO_w[3]) );
  AOI2BB2X1 U264 ( .B0(N240), .B1(n67), .A0N(n188), .A1N(n4), .Y(n20) );
  OAI221XL U265 ( .A0(n188), .A1(n11), .B0(n285), .B1(n12), .C0(n23), .Y(
        LO_w[2]) );
  AOI2BB2X1 U266 ( .B0(N239), .B1(n6), .A0N(n189), .A1N(n4), .Y(n23) );
  OAI221XL U267 ( .A0(n149), .A1(n14), .B0(n10), .B1(n207), .C0(n53), .Y(
        HI_w[9]) );
  OA22X1 U268 ( .A0(n56), .A1(n150), .B0(n208), .B1(n52), .Y(n53) );
  OAI221XL U269 ( .A0(n150), .A1(n36), .B0(n208), .B1(n5), .C0(n55), .Y(
        HI_w[8]) );
  OA22X1 U270 ( .A0(n58), .A1(n151), .B0(n209), .B1(n54), .Y(n55) );
  OAI221XL U271 ( .A0(n151), .A1(n36), .B0(n10), .B1(n209), .C0(n57), .Y(
        HI_w[7]) );
  OA22X1 U272 ( .A0(n56), .A1(n152), .B0(n210), .B1(n54), .Y(n57) );
  NOR2BX1 U273 ( .AN(N204), .B(n81), .Y(divisor_p[31]) );
  AO22X1 U274 ( .A0(n81), .A1(divisor[1]), .B0(N174), .B1(n87), .Y(
        divisor_p[1]) );
  AO22X1 U275 ( .A0(n83), .A1(divisor[2]), .B0(N175), .B1(n85), .Y(
        divisor_p[2]) );
  AO22X1 U276 ( .A0(n83), .A1(divisor[3]), .B0(N176), .B1(n85), .Y(
        divisor_p[3]) );
  AO22X1 U277 ( .A0(n83), .A1(divisor[4]), .B0(N177), .B1(n85), .Y(
        divisor_p[4]) );
  AO22X1 U278 ( .A0(n83), .A1(divisor[5]), .B0(N178), .B1(n85), .Y(
        divisor_p[5]) );
  AO22X1 U279 ( .A0(n83), .A1(divisor[6]), .B0(N179), .B1(n85), .Y(
        divisor_p[6]) );
  AO22X1 U280 ( .A0(n83), .A1(divisor[7]), .B0(N180), .B1(n85), .Y(
        divisor_p[7]) );
  AO22X1 U281 ( .A0(n83), .A1(divisor[8]), .B0(N181), .B1(n85), .Y(
        divisor_p[8]) );
  AO22X1 U282 ( .A0(n81), .A1(divisor[9]), .B0(N182), .B1(n85), .Y(
        divisor_p[9]) );
  AO22X1 U283 ( .A0(n81), .A1(divisor[10]), .B0(N183), .B1(n87), .Y(
        divisor_p[10]) );
  AO22X1 U284 ( .A0(n81), .A1(divisor[11]), .B0(N184), .B1(n87), .Y(
        divisor_p[11]) );
  AO22X1 U285 ( .A0(n81), .A1(divisor[12]), .B0(N185), .B1(n87), .Y(
        divisor_p[12]) );
  AO22X1 U286 ( .A0(n81), .A1(divisor[13]), .B0(N186), .B1(n87), .Y(
        divisor_p[13]) );
  AO22X1 U287 ( .A0(n81), .A1(divisor[14]), .B0(N187), .B1(n87), .Y(
        divisor_p[14]) );
  AO22X1 U288 ( .A0(n81), .A1(divisor[15]), .B0(N188), .B1(n85), .Y(
        divisor_p[15]) );
  AO22X1 U289 ( .A0(n81), .A1(divisor[16]), .B0(N189), .B1(n85), .Y(
        divisor_p[16]) );
  AO22X1 U290 ( .A0(n81), .A1(divisor[17]), .B0(N190), .B1(n87), .Y(
        divisor_p[17]) );
  AO22X1 U291 ( .A0(n81), .A1(divisor[18]), .B0(N191), .B1(n87), .Y(
        divisor_p[18]) );
  AO22X1 U292 ( .A0(n81), .A1(divisor[19]), .B0(N192), .B1(n87), .Y(
        divisor_p[19]) );
  AO22X1 U293 ( .A0(n81), .A1(divisor[20]), .B0(N193), .B1(n85), .Y(
        divisor_p[20]) );
  AO22X1 U294 ( .A0(n81), .A1(divisor[21]), .B0(N194), .B1(n85), .Y(
        divisor_p[21]) );
  AO22X1 U295 ( .A0(n81), .A1(divisor[22]), .B0(N195), .B1(n85), .Y(
        divisor_p[22]) );
  AO22X1 U296 ( .A0(n83), .A1(divisor[23]), .B0(N196), .B1(n85), .Y(
        divisor_p[23]) );
  AO22X1 U297 ( .A0(n83), .A1(divisor[24]), .B0(N197), .B1(n85), .Y(
        divisor_p[24]) );
  AO22X1 U298 ( .A0(n83), .A1(divisor[25]), .B0(N198), .B1(n85), .Y(
        divisor_p[25]) );
  AO22X1 U299 ( .A0(n83), .A1(divisor[26]), .B0(N199), .B1(n85), .Y(
        divisor_p[26]) );
  AO22X1 U300 ( .A0(n83), .A1(divisor[27]), .B0(N200), .B1(n85), .Y(
        divisor_p[27]) );
  AO22X1 U301 ( .A0(n83), .A1(divisor[28]), .B0(N201), .B1(n85), .Y(
        divisor_p[28]) );
  AO22X1 U302 ( .A0(n83), .A1(divisor[29]), .B0(N202), .B1(n85), .Y(
        divisor_p[29]) );
  AO22X1 U303 ( .A0(n83), .A1(divisor[30]), .B0(N203), .B1(n85), .Y(
        divisor_p[30]) );
  OAI2BB2XL U304 ( .B0(n159), .B1(n69), .A0N(N139), .A1N(n71), .Y(next_LO[31])
         );
  OAI2BB2XL U305 ( .B0(n160), .B1(n69), .A0N(N138), .A1N(n71), .Y(next_LO[30])
         );
  OAI2BB2XL U306 ( .B0(n161), .B1(n69), .A0N(N137), .A1N(n71), .Y(next_LO[29])
         );
  OAI2BB2XL U307 ( .B0(n162), .B1(n71), .A0N(N136), .A1N(n71), .Y(next_LO[28])
         );
  OAI2BB2XL U308 ( .B0(n163), .B1(n71), .A0N(N135), .A1N(n71), .Y(next_LO[27])
         );
  OAI2BB2XL U309 ( .B0(n164), .B1(n71), .A0N(N134), .A1N(n71), .Y(next_LO[26])
         );
  OAI2BB2XL U310 ( .B0(n165), .B1(n69), .A0N(N133), .A1N(n71), .Y(next_LO[25])
         );
  OAI2BB2XL U311 ( .B0(n166), .B1(n69), .A0N(N132), .A1N(n73), .Y(next_LO[24])
         );
  OAI2BB2XL U312 ( .B0(n167), .B1(n69), .A0N(N131), .A1N(n71), .Y(next_LO[23])
         );
  OAI2BB2XL U313 ( .B0(n75), .B1(n127), .A0N(N73), .A1N(n79), .Y(next_HI[31])
         );
  OAI2BB2XL U314 ( .B0(n77), .B1(n128), .A0N(N72), .A1N(n79), .Y(next_HI[30])
         );
  OAI2BB2XL U315 ( .B0(n75), .B1(n129), .A0N(N71), .A1N(n77), .Y(next_HI[29])
         );
  OAI2BB2XL U316 ( .B0(n75), .B1(n130), .A0N(N70), .A1N(n77), .Y(next_HI[28])
         );
  OAI2BB2XL U317 ( .B0(n75), .B1(n131), .A0N(N69), .A1N(n77), .Y(next_HI[27])
         );
  OAI2BB2XL U318 ( .B0(n75), .B1(n132), .A0N(N68), .A1N(n75), .Y(next_HI[26])
         );
  OAI2BB2XL U319 ( .B0(n75), .B1(n133), .A0N(N67), .A1N(n79), .Y(next_HI[25])
         );
  OAI2BB2XL U320 ( .B0(n75), .B1(n134), .A0N(N66), .A1N(n77), .Y(next_HI[24])
         );
  OAI2BB2XL U321 ( .B0(n75), .B1(n135), .A0N(N65), .A1N(n77), .Y(next_HI[23])
         );
  OAI2BB2XL U322 ( .B0(n75), .B1(n136), .A0N(N64), .A1N(n79), .Y(next_HI[22])
         );
  NOR2X1 U323 ( .A(state_r), .B(n219), .Y(div_stall) );
  CLKINVX1 U324 ( .A(div), .Y(n219) );
  OAI2BB2XL U325 ( .B0(n168), .B1(n69), .A0N(N130), .A1N(n71), .Y(next_LO[22])
         );
  OAI2BB2XL U326 ( .B0(n169), .B1(n69), .A0N(N129), .A1N(n73), .Y(next_LO[21])
         );
  OAI2BB2XL U327 ( .B0(n170), .B1(n69), .A0N(N128), .A1N(n71), .Y(next_LO[20])
         );
  OAI2BB2XL U328 ( .B0(n171), .B1(n69), .A0N(N127), .A1N(n73), .Y(next_LO[19])
         );
  OAI2BB2XL U329 ( .B0(n172), .B1(n69), .A0N(N126), .A1N(n73), .Y(next_LO[18])
         );
  OAI2BB2XL U330 ( .B0(n173), .B1(n69), .A0N(N125), .A1N(n73), .Y(next_LO[17])
         );
  OAI2BB2XL U331 ( .B0(n174), .B1(n69), .A0N(N124), .A1N(n73), .Y(next_LO[16])
         );
  OAI2BB2XL U332 ( .B0(n175), .B1(n69), .A0N(N123), .A1N(n73), .Y(next_LO[15])
         );
  OAI2BB2XL U333 ( .B0(n176), .B1(n69), .A0N(N122), .A1N(n73), .Y(next_LO[14])
         );
  OAI2BB2XL U334 ( .B0(n177), .B1(n69), .A0N(N121), .A1N(n73), .Y(next_LO[13])
         );
  CLKINVX1 U335 ( .A(diff[0]), .Y(n216) );
  OAI2BB2XL U336 ( .B0(n75), .B1(n137), .A0N(N63), .A1N(n79), .Y(next_HI[21])
         );
  OAI2BB2XL U337 ( .B0(n75), .B1(n138), .A0N(N62), .A1N(n79), .Y(next_HI[20])
         );
  OAI2BB2XL U338 ( .B0(n79), .B1(n139), .A0N(N61), .A1N(n79), .Y(next_HI[19])
         );
  OAI2BB2XL U339 ( .B0(n79), .B1(n140), .A0N(N60), .A1N(n79), .Y(next_HI[18])
         );
  OAI2BB2XL U340 ( .B0(n77), .B1(n141), .A0N(N59), .A1N(n79), .Y(next_HI[17])
         );
  OAI2BB2XL U341 ( .B0(sign_r[1]), .B1(n142), .A0N(N58), .A1N(n79), .Y(
        next_HI[16]) );
  OAI2BB2XL U342 ( .B0(n77), .B1(n143), .A0N(N57), .A1N(n79), .Y(next_HI[15])
         );
  OAI2BB2XL U343 ( .B0(sign_r[1]), .B1(n144), .A0N(N56), .A1N(n79), .Y(
        next_HI[14]) );
  OAI2BB2XL U344 ( .B0(sign_r[1]), .B1(n145), .A0N(N55), .A1N(n79), .Y(
        next_HI[13]) );
  OAI2BB2XL U345 ( .B0(sign_r[1]), .B1(n146), .A0N(N54), .A1N(n79), .Y(
        next_HI[12]) );
  AO22X1 U346 ( .A0(div_iter_r[5]), .A1(n85), .B0(n126), .B1(sign_r[0]), .Y(
        n124) );
  AO21X1 U347 ( .A0(n126), .A1(n75), .B0(n67), .Y(n125) );
  OAI2BB2XL U348 ( .B0(n183), .B1(n71), .A0N(N115), .A1N(n73), .Y(next_LO[7])
         );
  OAI2BB2XL U349 ( .B0(n184), .B1(n71), .A0N(N114), .A1N(n73), .Y(next_LO[6])
         );
  NOR4X1 U350 ( .A(n122), .B(n121), .C(n117), .D(n120), .Y(n116) );
  OR2X1 U351 ( .A(N273), .B(n119), .Y(n117) );
  OAI2BB2XL U352 ( .B0(n77), .B1(n147), .A0N(N53), .A1N(n75), .Y(next_HI[11])
         );
  OAI2BB2XL U353 ( .B0(n75), .B1(n148), .A0N(N52), .A1N(n75), .Y(next_HI[10])
         );
  OAI2BB2XL U354 ( .B0(n77), .B1(n149), .A0N(N51), .A1N(n75), .Y(next_HI[9])
         );
  OAI2BB2XL U355 ( .B0(n77), .B1(n150), .A0N(N50), .A1N(n75), .Y(next_HI[8])
         );
  OAI2BB2XL U356 ( .B0(n178), .B1(n69), .A0N(N120), .A1N(n73), .Y(next_LO[12])
         );
  OAI2BB2XL U357 ( .B0(n179), .B1(n69), .A0N(N119), .A1N(n73), .Y(next_LO[11])
         );
  CLKBUFX3 U358 ( .A(sign_r[1]), .Y(n77) );
  NAND2X1 U359 ( .A(n7), .B(n9), .Y(n259) );
  OAI21XL U360 ( .A0(N278), .A1(n219), .B0(n126), .Y(n9) );
  OAI2BB2XL U361 ( .B0(n77), .B1(n151), .A0N(N49), .A1N(n79), .Y(next_HI[7])
         );
  OAI2BB2XL U362 ( .B0(n77), .B1(n152), .A0N(N48), .A1N(n79), .Y(next_HI[6])
         );
  OAI2BB2XL U363 ( .B0(n77), .B1(n153), .A0N(N47), .A1N(n79), .Y(next_HI[5])
         );
  OAI2BB2XL U364 ( .B0(n77), .B1(n154), .A0N(N46), .A1N(n79), .Y(next_HI[4])
         );
  OAI2BB2XL U365 ( .B0(n77), .B1(n155), .A0N(N45), .A1N(n79), .Y(next_HI[3])
         );
  OAI2BB2XL U366 ( .B0(n75), .B1(n156), .A0N(N44), .A1N(n77), .Y(next_HI[2])
         );
  OAI2BB2XL U367 ( .B0(n77), .B1(n157), .A0N(N43), .A1N(n79), .Y(next_HI[1])
         );
  OAI2BB2XL U368 ( .B0(n75), .B1(n158), .A0N(N42), .A1N(n75), .Y(next_HI[0])
         );
  OAI2BB2XL U369 ( .B0(n180), .B1(n69), .A0N(N118), .A1N(n73), .Y(next_LO[10])
         );
  OAI2BB2XL U370 ( .B0(n181), .B1(n71), .A0N(N117), .A1N(n71), .Y(next_LO[9])
         );
  OAI2BB2XL U371 ( .B0(n182), .B1(n71), .A0N(N116), .A1N(n73), .Y(next_LO[8])
         );
  OAI2BB2XL U372 ( .B0(n185), .B1(n3), .A0N(N113), .A1N(n73), .Y(next_LO[5])
         );
  OAI2BB2XL U373 ( .B0(n186), .B1(n71), .A0N(N112), .A1N(n73), .Y(next_LO[4])
         );
  OAI2BB2XL U374 ( .B0(n187), .B1(n71), .A0N(N111), .A1N(n73), .Y(next_LO[3])
         );
  OAI2BB2XL U375 ( .B0(n188), .B1(n73), .A0N(N110), .A1N(n71), .Y(next_LO[2])
         );
  OAI2BB2XL U376 ( .B0(n189), .B1(n69), .A0N(N109), .A1N(n73), .Y(next_LO[1])
         );
  OAI2BB2XL U377 ( .B0(n69), .B1(n190), .A0N(N108), .A1N(n73), .Y(next_LO[0])
         );
  OAI2BB2XL U378 ( .B0(n119), .B1(n7), .A0N(N277), .A1N(n8), .Y(n258) );
  OAI2BB2XL U379 ( .B0(n120), .B1(n7), .A0N(N276), .A1N(n8), .Y(n257) );
  OAI2BB2XL U380 ( .B0(n121), .B1(n7), .A0N(N275), .A1N(n8), .Y(n256) );
  OAI2BB2XL U381 ( .B0(n122), .B1(n7), .A0N(N274), .A1N(n8), .Y(n255) );
  OAI2BB2XL U382 ( .B0(N273), .B1(n7), .A0N(N273), .A1N(n8), .Y(n260) );
  XOR2X1 U383 ( .A(\add_130/carry[5] ), .B(div_iter_r[5]), .Y(N278) );
endmodule


module Forwarding ( IDEX_RegRt, IDEX_RegRs, EXMEM_RegRd, MEMWB_RegRd, 
        EXMEM_RegWrite, MEMWB_RegWrite, forwardA, forwardB );
  input [4:0] IDEX_RegRt;
  input [4:0] IDEX_RegRs;
  input [4:0] EXMEM_RegRd;
  input [4:0] MEMWB_RegRd;
  output [1:0] forwardA;
  output [1:0] forwardB;
  input EXMEM_RegWrite, MEMWB_RegWrite;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n1, n2, n3, n4;

  NOR4X1 U1 ( .A(MEMWB_RegRd[0]), .B(MEMWB_RegRd[1]), .C(n22), .D(
        MEMWB_RegRd[2]), .Y(n7) );
  OR2XL U2 ( .A(MEMWB_RegRd[4]), .B(MEMWB_RegRd[3]), .Y(n22) );
  XNOR2X1 U3 ( .A(IDEX_RegRt[0]), .B(MEMWB_RegRd[0]), .Y(n16) );
  XNOR2X1 U4 ( .A(IDEX_RegRt[1]), .B(MEMWB_RegRd[1]), .Y(n18) );
  XNOR2X1 U5 ( .A(IDEX_RegRt[2]), .B(MEMWB_RegRd[2]), .Y(n17) );
  XNOR2X1 U6 ( .A(IDEX_RegRt[4]), .B(MEMWB_RegRd[4]), .Y(n15) );
  XNOR2X1 U7 ( .A(IDEX_RegRt[3]), .B(MEMWB_RegRd[3]), .Y(n19) );
  AND4X1 U8 ( .A(n8), .B(n9), .C(n10), .D(n11), .Y(forwardB[1]) );
  XOR2X1 U9 ( .A(n4), .B(IDEX_RegRt[1]), .Y(n8) );
  XOR2X1 U10 ( .A(n2), .B(IDEX_RegRt[0]), .Y(n9) );
  XOR2X1 U11 ( .A(n3), .B(IDEX_RegRt[2]), .Y(n10) );
  AND4X1 U12 ( .A(n2), .B(n4), .C(n29), .D(n3), .Y(n12) );
  NOR2X1 U13 ( .A(EXMEM_RegRd[4]), .B(EXMEM_RegRd[3]), .Y(n29) );
  NOR4X1 U14 ( .A(n12), .B(n1), .C(n13), .D(n14), .Y(n11) );
  XOR2X1 U15 ( .A(IDEX_RegRt[4]), .B(EXMEM_RegRd[4]), .Y(n13) );
  XOR2X1 U16 ( .A(IDEX_RegRt[3]), .B(EXMEM_RegRd[3]), .Y(n14) );
  NOR4X1 U17 ( .A(n5), .B(n6), .C(forwardB[1]), .D(n7), .Y(forwardB[0]) );
  NAND2X1 U18 ( .A(n15), .B(MEMWB_RegWrite), .Y(n6) );
  NAND4X1 U19 ( .A(n16), .B(n17), .C(n18), .D(n19), .Y(n5) );
  CLKINVX1 U20 ( .A(EXMEM_RegWrite), .Y(n1) );
  CLKINVX1 U21 ( .A(EXMEM_RegRd[1]), .Y(n4) );
  CLKINVX1 U22 ( .A(EXMEM_RegRd[2]), .Y(n3) );
  CLKINVX1 U23 ( .A(EXMEM_RegRd[0]), .Y(n2) );
  XNOR2X1 U24 ( .A(IDEX_RegRs[0]), .B(MEMWB_RegRd[0]), .Y(n31) );
  XNOR2X1 U25 ( .A(IDEX_RegRs[1]), .B(MEMWB_RegRd[1]), .Y(n33) );
  XNOR2X1 U26 ( .A(IDEX_RegRs[2]), .B(MEMWB_RegRd[2]), .Y(n32) );
  XNOR2X1 U27 ( .A(IDEX_RegRs[4]), .B(MEMWB_RegRd[4]), .Y(n30) );
  XNOR2X1 U28 ( .A(IDEX_RegRs[3]), .B(MEMWB_RegRd[3]), .Y(n34) );
  AND4X1 U29 ( .A(n23), .B(n24), .C(n25), .D(n26), .Y(forwardA[1]) );
  XOR2X1 U30 ( .A(n4), .B(IDEX_RegRs[1]), .Y(n23) );
  XOR2X1 U31 ( .A(n2), .B(IDEX_RegRs[0]), .Y(n24) );
  XOR2X1 U32 ( .A(n3), .B(IDEX_RegRs[2]), .Y(n25) );
  NOR4X1 U33 ( .A(n12), .B(n1), .C(n27), .D(n28), .Y(n26) );
  XOR2X1 U34 ( .A(IDEX_RegRs[3]), .B(EXMEM_RegRd[3]), .Y(n28) );
  XOR2X1 U35 ( .A(IDEX_RegRs[4]), .B(EXMEM_RegRd[4]), .Y(n27) );
  NOR4X1 U36 ( .A(n20), .B(n21), .C(forwardA[1]), .D(n7), .Y(forwardA[0]) );
  NAND2X1 U37 ( .A(n30), .B(MEMWB_RegWrite), .Y(n21) );
  NAND4X1 U38 ( .A(n31), .B(n32), .C(n33), .D(n34), .Y(n20) );
endmodule


module MIPS_Pipeline_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFXL U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFXL U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFXL U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFXL U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFXL U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  XOR3X1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  AND2X2 U1 ( .A(B[2]), .B(A[2]), .Y(n1) );
  XOR2X1 U2 ( .A(B[2]), .B(A[2]), .Y(SUM[2]) );
  CLKBUFX3 U3 ( .A(B[1]), .Y(SUM[1]) );
  CLKBUFX3 U4 ( .A(B[0]), .Y(SUM[0]) );
endmodule


module MIPS_Pipeline_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n16;
  wire   [31:1] carry;

  ADDFXL U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  AND2X2 U1 ( .A(B[2]), .B(A[2]), .Y(n1) );
  XOR2X1 U2 ( .A(A[30]), .B(n3), .Y(SUM[30]) );
  XOR2X1 U3 ( .A(A[29]), .B(n2), .Y(SUM[29]) );
  XOR2X1 U4 ( .A(A[28]), .B(n13), .Y(SUM[28]) );
  XOR2X1 U5 ( .A(A[27]), .B(n12), .Y(SUM[27]) );
  XOR2X1 U6 ( .A(A[26]), .B(n11), .Y(SUM[26]) );
  XOR2X1 U7 ( .A(A[25]), .B(n10), .Y(SUM[25]) );
  XOR2X1 U8 ( .A(A[24]), .B(n9), .Y(SUM[24]) );
  XNOR2X1 U9 ( .A(A[31]), .B(n16), .Y(SUM[31]) );
  NAND2X1 U10 ( .A(A[30]), .B(n3), .Y(n16) );
  AND2X2 U11 ( .A(A[28]), .B(n13), .Y(n2) );
  AND2X2 U12 ( .A(A[29]), .B(n2), .Y(n3) );
  AND2X2 U13 ( .A(A[18]), .B(carry[18]), .Y(n4) );
  AND2X2 U14 ( .A(A[19]), .B(n4), .Y(n5) );
  AND2X2 U15 ( .A(A[20]), .B(n5), .Y(n6) );
  AND2X2 U16 ( .A(A[21]), .B(n6), .Y(n7) );
  AND2X2 U17 ( .A(A[22]), .B(n7), .Y(n8) );
  AND2X2 U18 ( .A(A[23]), .B(n8), .Y(n9) );
  AND2X2 U19 ( .A(A[24]), .B(n9), .Y(n10) );
  AND2X2 U20 ( .A(A[25]), .B(n10), .Y(n11) );
  AND2X2 U21 ( .A(A[26]), .B(n11), .Y(n12) );
  AND2X2 U22 ( .A(A[27]), .B(n12), .Y(n13) );
  XOR2X1 U23 ( .A(A[18]), .B(carry[18]), .Y(SUM[18]) );
  XOR2X1 U24 ( .A(A[23]), .B(n8), .Y(SUM[23]) );
  XOR2X1 U25 ( .A(A[22]), .B(n7), .Y(SUM[22]) );
  XOR2X1 U26 ( .A(A[21]), .B(n6), .Y(SUM[21]) );
  XOR2X1 U27 ( .A(A[20]), .B(n5), .Y(SUM[20]) );
  XOR2X1 U28 ( .A(A[19]), .B(n4), .Y(SUM[19]) );
  XOR2X1 U29 ( .A(B[2]), .B(A[2]), .Y(SUM[2]) );
  CLKBUFX3 U30 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U31 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MIPS_Pipeline_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n30;

  XOR2X1 U1 ( .A(A[30]), .B(n27), .Y(SUM[30]) );
  XOR2X1 U2 ( .A(A[28]), .B(n25), .Y(SUM[28]) );
  XOR2X1 U3 ( .A(A[29]), .B(n26), .Y(SUM[29]) );
  XOR2X1 U4 ( .A(A[27]), .B(n24), .Y(SUM[27]) );
  XOR2X1 U5 ( .A(A[26]), .B(n23), .Y(SUM[26]) );
  XOR2X1 U6 ( .A(A[25]), .B(n22), .Y(SUM[25]) );
  XOR2X1 U7 ( .A(A[24]), .B(n21), .Y(SUM[24]) );
  XOR2X1 U8 ( .A(A[23]), .B(n20), .Y(SUM[23]) );
  XOR2X1 U9 ( .A(A[22]), .B(n19), .Y(SUM[22]) );
  XOR2X1 U10 ( .A(A[21]), .B(n18), .Y(SUM[21]) );
  XOR2X1 U11 ( .A(A[20]), .B(n17), .Y(SUM[20]) );
  XOR2X1 U12 ( .A(A[19]), .B(n16), .Y(SUM[19]) );
  XOR2X1 U13 ( .A(A[18]), .B(n15), .Y(SUM[18]) );
  XOR2X1 U14 ( .A(A[3]), .B(A[2]), .Y(SUM[3]) );
  XNOR2X1 U15 ( .A(A[31]), .B(n30), .Y(SUM[31]) );
  NAND2X1 U16 ( .A(A[30]), .B(n27), .Y(n30) );
  XOR2X1 U17 ( .A(A[6]), .B(n1), .Y(SUM[6]) );
  XOR2X1 U18 ( .A(A[5]), .B(n3), .Y(SUM[5]) );
  XOR2X1 U19 ( .A(A[4]), .B(n4), .Y(SUM[4]) );
  XOR2X1 U20 ( .A(A[17]), .B(n14), .Y(SUM[17]) );
  XOR2X1 U21 ( .A(A[16]), .B(n13), .Y(SUM[16]) );
  XOR2X1 U22 ( .A(A[15]), .B(n12), .Y(SUM[15]) );
  XOR2X1 U23 ( .A(A[14]), .B(n11), .Y(SUM[14]) );
  XOR2X1 U24 ( .A(A[13]), .B(n10), .Y(SUM[13]) );
  XOR2X1 U25 ( .A(A[12]), .B(n9), .Y(SUM[12]) );
  XOR2X1 U26 ( .A(A[11]), .B(n8), .Y(SUM[11]) );
  XOR2X1 U27 ( .A(A[10]), .B(n7), .Y(SUM[10]) );
  XOR2X1 U28 ( .A(A[9]), .B(n6), .Y(SUM[9]) );
  XOR2X1 U29 ( .A(A[8]), .B(n5), .Y(SUM[8]) );
  XOR2X1 U30 ( .A(A[7]), .B(n2), .Y(SUM[7]) );
  CLKINVX1 U31 ( .A(A[2]), .Y(SUM[2]) );
  AND2X2 U32 ( .A(A[5]), .B(n3), .Y(n1) );
  AND2X2 U33 ( .A(A[6]), .B(n1), .Y(n2) );
  AND2X2 U34 ( .A(A[4]), .B(n4), .Y(n3) );
  AND2X2 U35 ( .A(A[3]), .B(A[2]), .Y(n4) );
  AND2X2 U36 ( .A(A[7]), .B(n2), .Y(n5) );
  AND2X2 U37 ( .A(A[8]), .B(n5), .Y(n6) );
  AND2X2 U38 ( .A(A[9]), .B(n6), .Y(n7) );
  AND2X2 U39 ( .A(A[10]), .B(n7), .Y(n8) );
  AND2X2 U40 ( .A(A[11]), .B(n8), .Y(n9) );
  AND2X2 U41 ( .A(A[12]), .B(n9), .Y(n10) );
  AND2X2 U42 ( .A(A[13]), .B(n10), .Y(n11) );
  AND2X2 U43 ( .A(A[14]), .B(n11), .Y(n12) );
  AND2X2 U44 ( .A(A[15]), .B(n12), .Y(n13) );
  AND2X2 U45 ( .A(A[16]), .B(n13), .Y(n14) );
  AND2X2 U46 ( .A(A[17]), .B(n14), .Y(n15) );
  AND2X2 U47 ( .A(A[18]), .B(n15), .Y(n16) );
  AND2X2 U48 ( .A(A[19]), .B(n16), .Y(n17) );
  AND2X2 U49 ( .A(A[20]), .B(n17), .Y(n18) );
  AND2X2 U50 ( .A(A[21]), .B(n18), .Y(n19) );
  AND2X2 U51 ( .A(A[22]), .B(n19), .Y(n20) );
  AND2X2 U52 ( .A(A[23]), .B(n20), .Y(n21) );
  AND2X2 U53 ( .A(A[24]), .B(n21), .Y(n22) );
  AND2X2 U54 ( .A(A[25]), .B(n22), .Y(n23) );
  AND2X2 U55 ( .A(A[26]), .B(n23), .Y(n24) );
  AND2X2 U56 ( .A(A[27]), .B(n24), .Y(n25) );
  AND2X2 U57 ( .A(A[28]), .B(n25), .Y(n26) );
  AND2X2 U58 ( .A(A[29]), .B(n26), .Y(n27) );
  CLKBUFX3 U59 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U60 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MIPS_Pipeline ( i_clk, rst_n, ICACHE_ren, ICACHE_wen, ICACHE_addr, 
        ICACHE_wdata, ICACHE_stall, ICACHE_rdata, DCACHE_ren, DCACHE_wen, 
        DCACHE_addr, DCACHE_wdata, DCACHE_stall, DCACHE_rdata );
  output [29:0] ICACHE_addr;
  output [31:0] ICACHE_wdata;
  input [31:0] ICACHE_rdata;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input [31:0] DCACHE_rdata;
  input i_clk, rst_n, ICACHE_stall, DCACHE_stall;
  output ICACHE_ren, ICACHE_wen, DCACHE_ren, DCACHE_wen;
  wire   n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, inst_r_5, inst_r_4, inst_r_3, inst_r_2, inst_r_1,
         inst_r_0, PCSrc, IF_Flush, RegWrite, ALUSrc, RegDst, MemWrite,
         MemRead, MemtoReg, Jump, JumpR, raWrite, Branch, Shift, Mul, Div, HI,
         LO, taken, take, RegWrite_idex_r, RegWrite_exmem_r, RegWrite_memwb_r,
         stallJ, MemRead_idex_r, PCWrite, IFIDWrite, stall, Mul_idex_r,
         stall_mul, Div_idex_r, stall_div, take_r, N86, N87, N88, N89, N90,
         N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114,
         N115, N116, N117, take_w, RegWrite_idex_w, ALUSrc_idex_w,
         RegDst_idex_w, MemRead_idex_w, MemWrite_idex_w, MemtoReg_idex_w,
         Jump_idex_w, Shift_idex_w, Div_idex_w, Mul_idex_w, HI_idex_w,
         LO_idex_w, sign_ext_31, N298, N299, N300, N301, N302, N303, N304,
         N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315,
         N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326,
         N327, N328, N329, N346, n11, n13, n15, n29, n189, n221, n223, n253,
         n254, n257, n258, n259, n260, n262, n264, n266, n268, n270, n272,
         n274, n276, n278, n280, n282, n284, n286, n288, n290, n292, n294,
         n296, n298, n300, n302, n304, n306, n308, n310, n312, n314, n316,
         n318, n320, n322, n324, n326, n328, n330, n332, n334, n336, n338,
         n340, n342, n344, n346, n348, n350, n352, n354, n356, n358, n360,
         n362, n364, n366, n368, n370, n372, n374, n376, n378, n380, n382,
         n384, n386, n388, n390, n391, n393, n394, n395, n396, n399, n401,
         n403, n405, n407, n409, n411, n413, n415, n417, n419, n420, n422,
         n424, n426, n428, n430, n432, n434, n436, n438, n440, n442, n443,
         n445, n447, n449, n450, n452, n453, n455, n457, n459, n461, n463,
         n497, n498, n499, n500, n501, n502, n503, n504, n507, n508, n509,
         n510, n512, n513, n514, n515, n518, n519, n520, n521, n524, n525,
         n526, n527, n530, n531, n532, n533, n536, n537, n538, n539, n542,
         n543, n544, n545, n548, n549, n550, n551, n553, n554, n555, n557,
         n558, n559, n560, n563, n564, n565, n567, n568, n569, n570, n571,
         n574, n575, n576, n577, n580, n581, n582, n583, n586, n587, n588,
         n589, n592, n593, n594, n595, n598, n599, n600, n601, n604, n605,
         n606, n607, n610, n611, n612, n613, n616, n617, n618, n619, n622,
         n623, n625, n627, n628, n629, n630, n633, n634, n635, n636, n639,
         n640, n641, n642, n645, n646, n647, n648, n651, n652, n653, n654,
         n657, n658, n659, n660, n663, n664, n665, n666, n669, n670, n671,
         n672, n675, n676, n677, n678, n681, n682, n683, n684, n686, n687,
         n690, n691, n692, n693, n695, n696, n700, n701, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n790, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n947, n948, n949, n950, n951, n952, n954,
         n956, n958, n960, n962, n964, n966, n968, n970, n972, n974, n976,
         n978, n980, n982, n984, n986, n988, n990, n992, n994, n996, n998,
         n1000, n1002, n1004, n1006, n1008, n1010, n1012, n1014, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n75, n77, n79, n81, n83, n85, n87, n89, n91, n93,
         n95, n97, n99, n101, n103, n105, n107, n109, n111, n113, n115, n117,
         n119, n121, n123, n125, n127, n129, n131, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n183, n184, n185, n186, n187, n188, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n222, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n255, n256, n261, n263, n265, n267, n269, n271,
         n273, n275, n277, n279, n281, n283, n285, n287, n289, n291, n293,
         n295, n297, n299, n301, n303, n305, n307, n309, n311, n313, n315,
         n317, n319, n321, n323, n325, n327, n329, n331, n333, n335, n337,
         n339, n341, n343, n345, n347, n349, n351, n353, n355, n357, n359,
         n361, n363, n365, n367, n369, n371, n373, n375, n377, n379, n381,
         n383, n385, n387, n389, n392, n397, n398, n400, n402, n404, n406,
         n408, n410, n412, n414, n416, n418, n421, n423, n425, n427, n429,
         n431, n433, n435, n437, n439, n441, n444, n446, n448, n451, n454,
         n456, n458, n460, n462, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n505, n506, n511, n516, n517, n522, n523,
         n528, n529, n534, n535, n540, n541, n546, n547, n552, n556, n561,
         n562, n566, n572, n573, n578, n579, n584, n585, n590, n591, n596,
         n597, n602, n603, n608, n609, n614, n615, n620, n621, n624, n626,
         n631, n632, n637, n638, n643, n644, n649, n650, n655, n656, n661,
         n662, n667, n668, n673, n674, n679, n680, n685, n688, n689, n694,
         n697, n698, n699, n702, n703, n704, n705, n706, n707, n789, n791,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n953,
         n955, n957, n959, n961, n963, n965, n967, n969, n971, n973, n975,
         n977, n979, n981, n983, n985, n987, n989, n991, n993, n995, n997,
         n999, n1001, n1003, n1005, n1007, n1009, n1011, n1013, n1015, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683;
  wire   [1:0] PC_r;
  wire   [31:16] inst_r;
  wire   [1:0] ALUOp;
  wire   [4:0] RegRt_idex_r;
  wire   [4:0] RegRd_idex_r;
  wire   [5:0] Opcode_idex_r;
  wire   [4:0] RegRd_exmem_r;
  wire   [4:0] RegRd_memwb_r;
  wire   [1:0] ForwardJA;
  wire   [1:0] ForwardJB;
  wire   [31:0] Readdata1;
  wire   [31:0] Readdata2;
  wire   [5:0] Funct_idex_r;
  wire   [1:0] ALUOp_idex_r;
  wire   [3:0] ALUctrl;
  wire   [31:0] ALUin2;
  wire   [31:0] ALUresult;
  wire   [31:0] readreg1_forward;
  wire   [31:0] readreg2_forward;
  wire   [31:0] HI_mul;
  wire   [31:0] LO_mul;
  wire   [31:0] HI_div;
  wire   [31:0] LO_div;
  wire   [4:0] RegRs_idex_r;
  wire   [1:0] forwardA;
  wire   [1:0] forwardB;
  wire   [31:0] PC_4;
  wire   [31:0] PC_w;
  wire   [31:0] PC_4_r;
  wire   [31:0] PC_4_w;
  wire   [31:0] inst_w;
  wire   [1:0] ALUOp_idex_w;
  wire   [31:0] PC_4_idex_w;
  wire   [5:0] Opcode_idex_w;
  wire   [5:0] Funct_idex_w;
  wire   [4:0] RegRs_idex_w;
  wire   [4:0] RegRt_idex_w;
  wire   [4:0] RegRd_idex_w;
  wire   [4:0] shamt_idex_w;
  wire   [4:0] shamt_idex_r;
  wire   [31:0] readreg1_w;
  wire   [31:0] readreg2_w;
  wire   [31:0] sign_ext_w;
  wire   [14:6] sign_ext;
  assign ICACHE_wdata[0] = 1'b0;
  assign ICACHE_wdata[1] = 1'b0;
  assign ICACHE_wdata[2] = 1'b0;
  assign ICACHE_wdata[3] = 1'b0;
  assign ICACHE_wdata[4] = 1'b0;
  assign ICACHE_wdata[5] = 1'b0;
  assign ICACHE_wdata[6] = 1'b0;
  assign ICACHE_wdata[7] = 1'b0;
  assign ICACHE_wdata[8] = 1'b0;
  assign ICACHE_wdata[9] = 1'b0;
  assign ICACHE_wdata[10] = 1'b0;
  assign ICACHE_wdata[11] = 1'b0;
  assign ICACHE_wdata[12] = 1'b0;
  assign ICACHE_wdata[13] = 1'b0;
  assign ICACHE_wdata[14] = 1'b0;
  assign ICACHE_wdata[15] = 1'b0;
  assign ICACHE_wdata[16] = 1'b0;
  assign ICACHE_wdata[17] = 1'b0;
  assign ICACHE_wdata[18] = 1'b0;
  assign ICACHE_wdata[19] = 1'b0;
  assign ICACHE_wdata[20] = 1'b0;
  assign ICACHE_wdata[21] = 1'b0;
  assign ICACHE_wdata[22] = 1'b0;
  assign ICACHE_wdata[23] = 1'b0;
  assign ICACHE_wdata[24] = 1'b0;
  assign ICACHE_wdata[25] = 1'b0;
  assign ICACHE_wdata[26] = 1'b0;
  assign ICACHE_wdata[27] = 1'b0;
  assign ICACHE_wdata[28] = 1'b0;
  assign ICACHE_wdata[29] = 1'b0;
  assign ICACHE_wdata[30] = 1'b0;
  assign ICACHE_wdata[31] = 1'b0;
  assign ICACHE_wen = 1'b0;
  assign ICACHE_ren = 1'b1;

  OAI22X4 U1225 ( .A0(n1389), .A1(n1540), .B0(n1514), .B1(n205), .Y(ALUin2[9])
         );
  OAI22X4 U1231 ( .A0(n204), .A1(n1542), .B0(n1516), .B1(n206), .Y(ALUin2[8])
         );
  OAI22X4 U1237 ( .A0(n204), .A1(n1544), .B0(n1518), .B1(n207), .Y(ALUin2[7])
         );
  OAI22X4 U1261 ( .A0(n203), .A1(n1549), .B0(n1526), .B1(n205), .Y(ALUin2[3])
         );
  OAI22X4 U1285 ( .A0(n204), .A1(n1555), .B0(n1474), .B1(n207), .Y(ALUin2[29])
         );
  OAI22X4 U1291 ( .A0(n204), .A1(n1556), .B0(n1476), .B1(n205), .Y(ALUin2[28])
         );
  OAI22X4 U1297 ( .A0(n204), .A1(n1557), .B0(n1478), .B1(n205), .Y(ALUin2[27])
         );
  OAI22X4 U1309 ( .A0(n204), .A1(n1559), .B0(n1482), .B1(n44), .Y(ALUin2[25])
         );
  OAI22X4 U1321 ( .A0(n204), .A1(n1561), .B0(n1486), .B1(n205), .Y(ALUin2[23])
         );
  OAI22X4 U1333 ( .A0(n204), .A1(n1563), .B0(n1490), .B1(n205), .Y(ALUin2[21])
         );
  OAI22X4 U1345 ( .A0(n203), .A1(n1552), .B0(n1530), .B1(n206), .Y(ALUin2[1])
         );
  OAI22X4 U1351 ( .A0(n203), .A1(n1565), .B0(n1494), .B1(n206), .Y(ALUin2[19])
         );
  OAI22X4 U1375 ( .A0(n203), .A1(n1569), .B0(n1502), .B1(n208), .Y(ALUin2[15])
         );
  OAI22X4 U1387 ( .A0(n203), .A1(n1573), .B0(n1506), .B1(n206), .Y(ALUin2[13])
         );
  OAI22X4 U1393 ( .A0(n203), .A1(n1575), .B0(n1508), .B1(n207), .Y(ALUin2[12])
         );
  OAI22X4 U1399 ( .A0(n203), .A1(n1537), .B0(n1510), .B1(n207), .Y(ALUin2[11])
         );
  OAI22X4 U1405 ( .A0(n203), .A1(n1577), .B0(n1512), .B1(n207), .Y(ALUin2[10])
         );
  Control zctrl ( .inst({n72, inst_r[30:26]}), .funct({inst_r_5, inst_r_4, 
        inst_r_3, inst_r_2, inst_r_1, inst_r_0}), .eq(N346), .PCSrc(PCSrc), 
        .IF_Flush(IF_Flush), .RegWrite(RegWrite), .ALURsc(ALUSrc), .ALUOp(
        ALUOp), .RegDst(RegDst), .MemWrite(MemWrite), .MemRead(MemRead), 
        .MemtoReg(MemtoReg), .Jump(Jump), .JumpR(JumpR), .raWrite(raWrite), 
        .Branch(Branch), .Shift(Shift), .Mul(Mul), .Div(Div), .HI(HI), .LO(LO)
         );
  BranchPrd zbranchprd ( .clk(i_clk), .rst(n458), .taken(taken), .take(take), 
        .Branch(Branch) );
  forward_jump zforwardjump ( .JumpR(JumpR), .Branch(Branch), .RegJump(
        inst_r[25:21]), .RegRt(inst_r[20:16]), .IDEX_Opcode(Opcode_idex_r), 
        .IDEX_RegWrite(RegWrite_idex_r), .IDEX_RegRt(RegRt_idex_r), 
        .IDEX_RegRd(RegRd_idex_r), .EXMEM_RegWrite(RegWrite_exmem_r), 
        .EXMEM_MemRead(DCACHE_ren), .EXMEM_RegRd(RegRd_exmem_r), 
        .MEMWB_RegWrite(RegWrite_memwb_r), .MEMWB_RegRd(RegRd_memwb_r), 
        .ForwardJA(ForwardJA), .ForwardJB(ForwardJB), .stallJ(stallJ) );
  HazardDetection zhd ( .opcode({n72, inst_r[30:26]}), .IDEX_MemRead(
        MemRead_idex_r), .IDEX_RegRt(RegRt_idex_r), .IFID_RegRs(inst_r[25:21]), 
        .IFID_RegRt(inst_r[20:16]), .PCWrite(PCWrite), .IFIDWrite(IFIDWrite), 
        .stall(stall) );
  register zregister ( .clk(i_clk), .rst_n(n458), .RegWrite(RegWrite_memwb_r), 
        .ReadReg1(inst_r[25:21]), .ReadReg2(inst_r[20:16]), .WriteReg({
        RegRd_memwb_r[4:2], n73, RegRd_memwb_r[0]}), .WriteData({n1430, n1431, 
        n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, 
        n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, 
        n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461}), 
        .ReadData1(Readdata1), .ReadData2(Readdata2) );
  aluCtrl zaluCtrl ( .opcode(Opcode_idex_r), .funct(Funct_idex_r), .ALUOp(
        ALUOp_idex_r), .ctrl(ALUctrl) );
  alu zalu ( .ctrl(ALUctrl), .x({n1370, n1369, n1367, n1366, n1365, n1364, 
        n1363, n1362, n1361, n1360, n1359, n1358, n1356, n1355, n1354, n1353, 
        n1352, n1351, n1350, n1349, n1348, n1347, n1377, n1376, n1375, n1374, 
        n1373, n1372, n1371, n1368, n1357, n1346}), .y(ALUin2), .out(ALUresult) );
  mul zmul ( .clk(i_clk), .rst(n458), .mul(Mul_idex_r), .multiplicand(
        readreg1_forward), .LO({n454, readreg2_forward[30:0]}), .next_HI(
        HI_mul), .next_LO(LO_mul), .mul_stall(stall_mul) );
  div zdiv ( .clk(i_clk), .rst(n458), .div(Div_idex_r), .divisor({n454, 
        readreg2_forward[30:0]}), .LO(readreg1_forward), .next_HI(HI_div), 
        .next_LO(LO_div), .div_stall(stall_div) );
  Forwarding zforwarding ( .IDEX_RegRt(RegRt_idex_r), .IDEX_RegRs(RegRs_idex_r), .EXMEM_RegRd(RegRd_exmem_r), .MEMWB_RegRd({RegRd_memwb_r[4], n70, n71, 
        RegRd_memwb_r[1:0]}), .EXMEM_RegWrite(RegWrite_exmem_r), 
        .MEMWB_RegWrite(RegWrite_memwb_r), .forwardA(forwardA), .forwardB(
        forwardB) );
  MIPS_Pipeline_DW01_add_0 add_297 ( .A({n198, n198, n198, n198, n198, n198, 
        n198, n198, n198, n198, n198, n198, n198, n198, n198, sign_ext, 
        inst_r_5, inst_r_4, inst_r_3, inst_r_2, inst_r_1, inst_r_0, 1'b0, 1'b0}), .B(PC_4_r), .CI(1'b0), .SUM({N329, N328, N327, N326, N325, N324, N323, N322, 
        N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, 
        N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298}) );
  MIPS_Pipeline_DW01_add_1 add_188 ( .A(PC_4), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        ICACHE_rdata[15:0], 1'b0, 1'b0}), .CI(1'b0), .SUM({N117, N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86}) );
  MIPS_Pipeline_DW01_add_2 add_174 ( .A({ICACHE_addr, PC_r}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(PC_4) );
  DFFRX1 \PC_4_r_reg[0]  ( .D(PC_4_w[0]), .CK(i_clk), .RN(n460), .Q(PC_4_r[0]), 
        .QN(n1383) );
  DFFRX1 \PC_4_r_reg[1]  ( .D(PC_4_w[1]), .CK(i_clk), .RN(n460), .Q(PC_4_r[1]), 
        .QN(n1382) );
  DFFRX1 \PC_4_idex_r_reg[0]  ( .D(PC_4_idex_w[0]), .CK(i_clk), .RN(n460), 
        .QN(n1101) );
  DFFRX1 \PC_4_idex_r_reg[1]  ( .D(PC_4_idex_w[1]), .CK(i_clk), .RN(n460), 
        .QN(n1076) );
  DFFRX1 \PC_4_idex_r_reg[2]  ( .D(PC_4_idex_w[2]), .CK(i_clk), .RN(n460), 
        .QN(n1074) );
  DFFRX1 \PC_4_idex_r_reg[3]  ( .D(PC_4_idex_w[3]), .CK(i_clk), .RN(n462), 
        .QN(n1072) );
  DFFRX1 \PC_4_idex_r_reg[4]  ( .D(PC_4_idex_w[4]), .CK(i_clk), .RN(n462), 
        .QN(n1070) );
  DFFRX1 \PC_4_idex_r_reg[5]  ( .D(PC_4_idex_w[5]), .CK(i_clk), .RN(n462), 
        .QN(n1068) );
  DFFRX1 \PC_4_idex_r_reg[6]  ( .D(PC_4_idex_w[6]), .CK(i_clk), .RN(n462), 
        .QN(n1066) );
  DFFRX1 \PC_4_idex_r_reg[7]  ( .D(PC_4_idex_w[7]), .CK(i_clk), .RN(n462), 
        .QN(n1064) );
  DFFRX1 \PC_4_idex_r_reg[8]  ( .D(PC_4_idex_w[8]), .CK(i_clk), .RN(n462), 
        .QN(n1062) );
  DFFRX1 \PC_4_idex_r_reg[9]  ( .D(PC_4_idex_w[9]), .CK(i_clk), .RN(n462), 
        .QN(n1060) );
  DFFRX1 \PC_4_idex_r_reg[10]  ( .D(PC_4_idex_w[10]), .CK(i_clk), .RN(n462), 
        .QN(n1058) );
  DFFRX1 \PC_4_idex_r_reg[11]  ( .D(PC_4_idex_w[11]), .CK(i_clk), .RN(n462), 
        .QN(n1056) );
  DFFRX1 \PC_4_idex_r_reg[12]  ( .D(PC_4_idex_w[12]), .CK(i_clk), .RN(n464), 
        .QN(n1054) );
  DFFRX1 \PC_4_idex_r_reg[13]  ( .D(PC_4_idex_w[13]), .CK(i_clk), .RN(n464), 
        .QN(n1052) );
  DFFRX1 \PC_4_idex_r_reg[14]  ( .D(PC_4_idex_w[14]), .CK(i_clk), .RN(n464), 
        .QN(n1050) );
  DFFRX1 \PC_4_idex_r_reg[15]  ( .D(PC_4_idex_w[15]), .CK(i_clk), .RN(n464), 
        .QN(n1048) );
  DFFRX1 \PC_4_idex_r_reg[16]  ( .D(PC_4_idex_w[16]), .CK(i_clk), .RN(n464), 
        .QN(n1046) );
  DFFRX1 \PC_4_idex_r_reg[17]  ( .D(PC_4_idex_w[17]), .CK(i_clk), .RN(n464), 
        .QN(n1044) );
  DFFRX1 \PC_4_idex_r_reg[18]  ( .D(PC_4_idex_w[18]), .CK(i_clk), .RN(n464), 
        .QN(n1042) );
  DFFRX1 \PC_4_idex_r_reg[19]  ( .D(PC_4_idex_w[19]), .CK(i_clk), .RN(n464), 
        .QN(n1040) );
  DFFRX1 \PC_4_idex_r_reg[20]  ( .D(PC_4_idex_w[20]), .CK(i_clk), .RN(n465), 
        .QN(n1038) );
  DFFRX1 \PC_4_idex_r_reg[21]  ( .D(PC_4_idex_w[21]), .CK(i_clk), .RN(n471), 
        .QN(n1036) );
  DFFRX1 \PC_4_idex_r_reg[22]  ( .D(PC_4_idex_w[22]), .CK(i_clk), .RN(n472), 
        .QN(n1034) );
  DFFRX1 \PC_4_idex_r_reg[23]  ( .D(PC_4_idex_w[23]), .CK(i_clk), .RN(n472), 
        .QN(n1032) );
  DFFRX1 \PC_4_idex_r_reg[24]  ( .D(PC_4_idex_w[24]), .CK(i_clk), .RN(n472), 
        .QN(n1030) );
  DFFRX1 \PC_4_idex_r_reg[25]  ( .D(PC_4_idex_w[25]), .CK(i_clk), .RN(n472), 
        .QN(n1028) );
  DFFRX1 \PC_4_idex_r_reg[26]  ( .D(PC_4_idex_w[26]), .CK(i_clk), .RN(n472), 
        .QN(n1026) );
  DFFRX1 \PC_4_idex_r_reg[27]  ( .D(PC_4_idex_w[27]), .CK(i_clk), .RN(n472), 
        .QN(n1024) );
  DFFRX1 \PC_4_idex_r_reg[28]  ( .D(PC_4_idex_w[28]), .CK(i_clk), .RN(n472), 
        .QN(n1022) );
  DFFRX1 \PC_4_idex_r_reg[29]  ( .D(PC_4_idex_w[29]), .CK(i_clk), .RN(n472), 
        .QN(n1020) );
  DFFRX1 \PC_4_idex_r_reg[30]  ( .D(PC_4_idex_w[30]), .CK(i_clk), .RN(n472), 
        .QN(n1018) );
  DFFRX1 \PC_4_idex_r_reg[31]  ( .D(PC_4_idex_w[31]), .CK(i_clk), .RN(n469), 
        .QN(n1103) );
  DFFRX1 \PC_4_r_reg[30]  ( .D(PC_4_w[30]), .CK(i_clk), .RN(n472), .Q(
        PC_4_r[30]), .QN(n1379) );
  DFFRX1 \PC_4_r_reg[31]  ( .D(PC_4_w[31]), .CK(i_clk), .RN(n468), .Q(
        PC_4_r[31]), .QN(n1378) );
  DFFRX1 MemtoReg_exmem_r_reg ( .D(n1244), .CK(i_clk), .RN(n466), .QN(n1104)
         );
  DFFRX1 MemtoReg_idex_r_reg ( .D(MemtoReg_idex_w), .CK(i_clk), .RN(n466), 
        .QN(n1099) );
  DFFRX1 MemWrite_idex_r_reg ( .D(MemWrite_idex_w), .CK(i_clk), .RN(n466), 
        .QN(n1095) );
  DFFRX1 Jump_idex_r_reg ( .D(Jump_idex_w), .CK(i_clk), .RN(n465), .QN(n1396)
         );
  DFFRX1 RegDst_idex_r_reg ( .D(RegDst_idex_w), .CK(i_clk), .RN(n466), .QN(
        n1090) );
  DFFRX1 RegWrite_idex_r_reg ( .D(RegWrite_idex_w), .CK(i_clk), .RN(n466), .Q(
        RegWrite_idex_r), .QN(n1093) );
  DFFRX1 \PC_4_r_reg[23]  ( .D(PC_4_w[23]), .CK(i_clk), .RN(n472), .Q(
        PC_4_r[23]), .QN(n885) );
  DFFRX1 \PC_4_r_reg[24]  ( .D(PC_4_w[24]), .CK(i_clk), .RN(n472), .Q(
        PC_4_r[24]), .QN(n886) );
  DFFRX1 \PC_4_r_reg[25]  ( .D(PC_4_w[25]), .CK(i_clk), .RN(n472), .Q(
        PC_4_r[25]), .QN(n887) );
  DFFRX1 \PC_4_r_reg[26]  ( .D(PC_4_w[26]), .CK(i_clk), .RN(n472), .Q(
        PC_4_r[26]), .QN(n888) );
  DFFRX1 \PC_4_r_reg[27]  ( .D(PC_4_w[27]), .CK(i_clk), .RN(n472), .Q(
        PC_4_r[27]), .QN(n889) );
  DFFRX1 \PC_4_r_reg[28]  ( .D(PC_4_w[28]), .CK(i_clk), .RN(n472), .Q(
        PC_4_r[28]), .QN(n1381) );
  DFFRX1 \PC_4_r_reg[29]  ( .D(PC_4_w[29]), .CK(i_clk), .RN(n472), .Q(
        PC_4_r[29]), .QN(n1380) );
  DFFRX1 MemRead_idex_r_reg ( .D(MemRead_idex_w), .CK(i_clk), .RN(n466), .Q(
        MemRead_idex_r), .QN(n1097) );
  DFFRX1 \Funct_idex_r_reg[3]  ( .D(Funct_idex_w[3]), .CK(i_clk), .RN(n467), 
        .Q(Funct_idex_r[3]), .QN(n796) );
  DFFRX1 \Funct_idex_r_reg[2]  ( .D(Funct_idex_w[2]), .CK(i_clk), .RN(n467), 
        .Q(Funct_idex_r[2]), .QN(n795) );
  DFFRX1 \Funct_idex_r_reg[1]  ( .D(Funct_idex_w[1]), .CK(i_clk), .RN(n468), 
        .Q(Funct_idex_r[1]), .QN(n794) );
  DFFRX1 \Funct_idex_r_reg[0]  ( .D(Funct_idex_w[0]), .CK(i_clk), .RN(n460), 
        .Q(Funct_idex_r[0]), .QN(n793) );
  DFFRX1 Div_idex_r_reg ( .D(Div_idex_w), .CK(i_clk), .RN(n469), .Q(Div_idex_r), .QN(n1397) );
  DFFRX1 \Funct_idex_r_reg[4]  ( .D(Funct_idex_w[4]), .CK(i_clk), .RN(n467), 
        .Q(Funct_idex_r[4]), .QN(n797) );
  DFFRX1 \Opcode_idex_r_reg[3]  ( .D(Opcode_idex_w[3]), .CK(i_clk), .RN(n467), 
        .Q(Opcode_idex_r[3]), .QN(n869) );
  DFFRX1 \Opcode_idex_r_reg[2]  ( .D(Opcode_idex_w[2]), .CK(i_clk), .RN(n467), 
        .Q(Opcode_idex_r[2]), .QN(n868) );
  DFFRX1 \RegRd_idex_r_reg[0]  ( .D(RegRd_idex_w[0]), .CK(i_clk), .RN(n466), 
        .Q(RegRd_idex_r[0]), .QN(n1089) );
  DFFRX1 \RegRd_idex_r_reg[2]  ( .D(RegRd_idex_w[2]), .CK(i_clk), .RN(n460), 
        .Q(RegRd_idex_r[2]), .QN(n1081) );
  DFFRX1 \HI_r_reg[20]  ( .D(n1003), .CK(i_clk), .RN(n471), .Q(n69), .QN(n812)
         );
  DFFRX1 \HI_r_reg[21]  ( .D(n1001), .CK(i_clk), .RN(n471), .Q(n68), .QN(n813)
         );
  DFFRX1 \HI_r_reg[22]  ( .D(n999), .CK(i_clk), .RN(n471), .Q(n67), .QN(n814)
         );
  DFFRX1 \HI_r_reg[23]  ( .D(n997), .CK(i_clk), .RN(n471), .Q(n66), .QN(n815)
         );
  DFFRX1 \HI_r_reg[24]  ( .D(n995), .CK(i_clk), .RN(n471), .Q(n65), .QN(n816)
         );
  DFFRX1 \HI_r_reg[25]  ( .D(n993), .CK(i_clk), .RN(n471), .Q(n64), .QN(n817)
         );
  DFFRX1 \HI_r_reg[26]  ( .D(n991), .CK(i_clk), .RN(n471), .Q(n63), .QN(n818)
         );
  DFFRX1 \HI_r_reg[27]  ( .D(n989), .CK(i_clk), .RN(n471), .Q(n62), .QN(n819)
         );
  DFFRX1 \HI_r_reg[28]  ( .D(n987), .CK(i_clk), .RN(n471), .Q(n61), .QN(n820)
         );
  DFFRX1 \HI_r_reg[29]  ( .D(n985), .CK(i_clk), .RN(n471), .Q(n60), .QN(n821)
         );
  DFFRX1 \HI_r_reg[30]  ( .D(n981), .CK(i_clk), .RN(n471), .Q(n59), .QN(n823)
         );
  DFFRX1 \HI_r_reg[31]  ( .D(n979), .CK(i_clk), .RN(n458), .Q(n58), .QN(n824)
         );
  DFFRX1 \LO_r_reg[20]  ( .D(n940), .CK(i_clk), .RN(n470), .Q(n57), .QN(n845)
         );
  DFFRX1 \LO_r_reg[21]  ( .D(n939), .CK(i_clk), .RN(n470), .Q(n56), .QN(n846)
         );
  DFFRX1 \LO_r_reg[22]  ( .D(n938), .CK(i_clk), .RN(n470), .Q(n55), .QN(n847)
         );
  DFFRX1 \LO_r_reg[23]  ( .D(n937), .CK(i_clk), .RN(n470), .Q(n54), .QN(n848)
         );
  DFFRX1 \LO_r_reg[24]  ( .D(n936), .CK(i_clk), .RN(n470), .Q(n53), .QN(n849)
         );
  DFFRX1 \LO_r_reg[25]  ( .D(n935), .CK(i_clk), .RN(n470), .Q(n52), .QN(n850)
         );
  DFFRX1 \LO_r_reg[26]  ( .D(n934), .CK(i_clk), .RN(n470), .Q(n51), .QN(n851)
         );
  DFFRX1 \LO_r_reg[27]  ( .D(n933), .CK(i_clk), .RN(n470), .Q(n50), .QN(n852)
         );
  DFFRX1 \LO_r_reg[28]  ( .D(n932), .CK(i_clk), .RN(n470), .Q(n49), .QN(n853)
         );
  DFFRX1 \LO_r_reg[29]  ( .D(n931), .CK(i_clk), .RN(n470), .Q(n48), .QN(n854)
         );
  DFFRX1 \LO_r_reg[30]  ( .D(n929), .CK(i_clk), .RN(n470), .Q(n47), .QN(n856)
         );
  DFFRX1 \LO_r_reg[31]  ( .D(n928), .CK(i_clk), .RN(n470), .Q(n46), .QN(n857)
         );
  DFFRX1 \PC_4_r_reg[15]  ( .D(PC_4_w[15]), .CK(i_clk), .RN(n464), .Q(
        PC_4_r[15]), .QN(n877) );
  DFFRX1 \PC_4_r_reg[16]  ( .D(PC_4_w[16]), .CK(i_clk), .RN(n464), .Q(
        PC_4_r[16]), .QN(n878) );
  DFFRX1 \PC_4_r_reg[17]  ( .D(PC_4_w[17]), .CK(i_clk), .RN(n464), .Q(
        PC_4_r[17]), .QN(n879) );
  DFFRX1 \PC_4_r_reg[18]  ( .D(PC_4_w[18]), .CK(i_clk), .RN(n464), .Q(
        PC_4_r[18]), .QN(n880) );
  DFFRX1 \PC_4_r_reg[19]  ( .D(PC_4_w[19]), .CK(i_clk), .RN(n464), .Q(
        PC_4_r[19]), .QN(n881) );
  DFFRX1 \PC_4_r_reg[20]  ( .D(PC_4_w[20]), .CK(i_clk), .RN(n464), .Q(
        PC_4_r[20]), .QN(n882) );
  DFFRX1 \PC_4_r_reg[21]  ( .D(PC_4_w[21]), .CK(i_clk), .RN(n471), .Q(
        PC_4_r[21]), .QN(n883) );
  DFFRX1 \PC_4_r_reg[22]  ( .D(PC_4_w[22]), .CK(i_clk), .RN(n472), .Q(
        PC_4_r[22]), .QN(n884) );
  DFFRX1 \RegRd_idex_r_reg[4]  ( .D(RegRd_idex_w[4]), .CK(i_clk), .RN(n460), 
        .Q(RegRd_idex_r[4]), .QN(n1395) );
  DFFRX1 \RegRd_idex_r_reg[3]  ( .D(RegRd_idex_w[3]), .CK(i_clk), .RN(n460), 
        .Q(RegRd_idex_r[3]), .QN(n1084) );
  DFFRX1 \RegRd_idex_r_reg[1]  ( .D(RegRd_idex_w[1]), .CK(i_clk), .RN(n460), 
        .Q(RegRd_idex_r[1]), .QN(n1078) );
  DFFRX1 \Opcode_idex_r_reg[4]  ( .D(Opcode_idex_w[4]), .CK(i_clk), .RN(n467), 
        .Q(Opcode_idex_r[4]), .QN(n870) );
  DFFRX1 \Opcode_idex_r_reg[1]  ( .D(Opcode_idex_w[1]), .CK(i_clk), .RN(n467), 
        .Q(Opcode_idex_r[1]), .QN(n867) );
  DFFRX1 \Opcode_idex_r_reg[0]  ( .D(Opcode_idex_w[0]), .CK(i_clk), .RN(n467), 
        .Q(Opcode_idex_r[0]), .QN(n866) );
  DFFRX1 Mul_idex_r_reg ( .D(Mul_idex_w), .CK(i_clk), .RN(n466), .Q(Mul_idex_r), .QN(n865) );
  DFFRX1 \inst_r_reg[28]  ( .D(inst_w[28]), .CK(i_clk), .RN(n467), .Q(
        inst_r[28]), .QN(n911) );
  DFFRX1 \Funct_idex_r_reg[5]  ( .D(Funct_idex_w[5]), .CK(i_clk), .RN(n467), 
        .Q(Funct_idex_r[5]), .QN(n798) );
  DFFRX1 \Opcode_idex_r_reg[5]  ( .D(Opcode_idex_w[5]), .CK(i_clk), .RN(n467), 
        .Q(Opcode_idex_r[5]), .QN(n871) );
  DFFRX1 \ALUresult2_r_reg[18]  ( .D(n1194), .CK(i_clk), .RN(n464), .QN(n1041)
         );
  DFFRX1 \ALUresult2_r_reg[19]  ( .D(n1192), .CK(i_clk), .RN(n464), .QN(n1039)
         );
  DFFRX1 \ALUresult2_r_reg[20]  ( .D(n1190), .CK(i_clk), .RN(n471), .QN(n1037)
         );
  DFFRX1 \ALUresult2_r_reg[21]  ( .D(n1188), .CK(i_clk), .RN(n472), .QN(n1035)
         );
  DFFRX1 \ALUresult2_r_reg[22]  ( .D(n1186), .CK(i_clk), .RN(n472), .QN(n1033)
         );
  DFFRX1 \ALUresult2_r_reg[23]  ( .D(n1184), .CK(i_clk), .RN(n472), .QN(n1031)
         );
  DFFRX1 \ALUresult2_r_reg[24]  ( .D(n1182), .CK(i_clk), .RN(n472), .QN(n1029)
         );
  DFFRX1 \ALUresult2_r_reg[25]  ( .D(n1180), .CK(i_clk), .RN(n472), .QN(n1027)
         );
  DFFRX1 \ALUresult2_r_reg[26]  ( .D(n1178), .CK(i_clk), .RN(n472), .QN(n1025)
         );
  DFFRX1 \ALUresult2_r_reg[27]  ( .D(n1176), .CK(i_clk), .RN(n472), .QN(n1023)
         );
  DFFRX1 \ALUresult2_r_reg[28]  ( .D(n1174), .CK(i_clk), .RN(n472), .QN(n1021)
         );
  DFFRX1 \ALUresult2_r_reg[29]  ( .D(n1172), .CK(i_clk), .RN(n472), .QN(n1019)
         );
  DFFRX1 \ALUresult2_r_reg[30]  ( .D(n1170), .CK(i_clk), .RN(n473), .QN(n1017)
         );
  DFFRX1 \PC_4_r_reg[7]  ( .D(PC_4_w[7]), .CK(i_clk), .RN(n462), .Q(PC_4_r[7]), 
        .QN(n895) );
  DFFRX1 \PC_4_r_reg[8]  ( .D(PC_4_w[8]), .CK(i_clk), .RN(n462), .Q(PC_4_r[8]), 
        .QN(n896) );
  DFFRX1 \PC_4_r_reg[9]  ( .D(PC_4_w[9]), .CK(i_clk), .RN(n462), .Q(PC_4_r[9]), 
        .QN(n897) );
  DFFRX1 \PC_4_r_reg[10]  ( .D(PC_4_w[10]), .CK(i_clk), .RN(n462), .Q(
        PC_4_r[10]), .QN(n872) );
  DFFRX1 \PC_4_r_reg[11]  ( .D(PC_4_w[11]), .CK(i_clk), .RN(n462), .Q(
        PC_4_r[11]), .QN(n873) );
  DFFRX1 \PC_4_r_reg[12]  ( .D(PC_4_w[12]), .CK(i_clk), .RN(n464), .Q(
        PC_4_r[12]), .QN(n874) );
  DFFRX1 \PC_4_r_reg[13]  ( .D(PC_4_w[13]), .CK(i_clk), .RN(n464), .Q(
        PC_4_r[13]), .QN(n875) );
  DFFRX1 \PC_4_r_reg[14]  ( .D(PC_4_w[14]), .CK(i_clk), .RN(n464), .Q(
        PC_4_r[14]), .QN(n876) );
  DFFRX1 \inst_r_reg[5]  ( .D(inst_w[5]), .CK(i_clk), .RN(n466), .Q(inst_r_5), 
        .QN(n952) );
  DFFRX1 MemRead_exmem_r_reg ( .D(n1243), .CK(i_clk), .RN(n466), .Q(DCACHE_ren), .QN(n1098) );
  DFFRX1 \ALUresult2_r_reg[11]  ( .D(n1208), .CK(i_clk), .RN(n464), .QN(n1055)
         );
  DFFRX1 \ALUresult2_r_reg[12]  ( .D(n1206), .CK(i_clk), .RN(n464), .QN(n1053)
         );
  DFFRX1 \ALUresult2_r_reg[13]  ( .D(n1204), .CK(i_clk), .RN(n464), .QN(n1051)
         );
  DFFRX1 \ALUresult2_r_reg[14]  ( .D(n1202), .CK(i_clk), .RN(n464), .QN(n1049)
         );
  DFFRX1 \ALUresult2_r_reg[15]  ( .D(n1200), .CK(i_clk), .RN(n464), .QN(n1047)
         );
  DFFRX1 \ALUresult2_r_reg[16]  ( .D(n1198), .CK(i_clk), .RN(n464), .QN(n1045)
         );
  DFFRX1 \ALUresult2_r_reg[17]  ( .D(n1196), .CK(i_clk), .RN(n464), .QN(n1043)
         );
  DFFRX1 \PC_4_r_reg[2]  ( .D(PC_4_w[2]), .CK(i_clk), .RN(n460), .Q(PC_4_r[2]), 
        .QN(n890) );
  DFFRX1 \PC_4_r_reg[3]  ( .D(PC_4_w[3]), .CK(i_clk), .RN(n462), .Q(PC_4_r[3]), 
        .QN(n891) );
  DFFRX1 \PC_4_r_reg[4]  ( .D(PC_4_w[4]), .CK(i_clk), .RN(n462), .Q(PC_4_r[4]), 
        .QN(n892) );
  DFFRX1 \PC_4_r_reg[5]  ( .D(PC_4_w[5]), .CK(i_clk), .RN(n462), .Q(PC_4_r[5]), 
        .QN(n893) );
  DFFRX1 \PC_4_r_reg[6]  ( .D(PC_4_w[6]), .CK(i_clk), .RN(n462), .Q(PC_4_r[6]), 
        .QN(n894) );
  DFFRX1 \inst_r_reg[2]  ( .D(inst_w[2]), .CK(i_clk), .RN(n467), .Q(inst_r_2), 
        .QN(n949) );
  DFFRX1 \inst_r_reg[0]  ( .D(inst_w[0]), .CK(i_clk), .RN(n460), .Q(inst_r_0), 
        .QN(n947) );
  DFFRX1 \inst_r_reg[25]  ( .D(inst_w[25]), .CK(i_clk), .RN(n467), .Q(
        inst_r[25]), .QN(n908) );
  DFFRX1 \inst_r_reg[24]  ( .D(inst_w[24]), .CK(i_clk), .RN(n467), .Q(
        inst_r[24]), .QN(n907) );
  DFFRX1 \inst_r_reg[4]  ( .D(inst_w[4]), .CK(i_clk), .RN(n467), .Q(inst_r_4), 
        .QN(n951) );
  DFFRX1 \inst_r_reg[23]  ( .D(inst_w[23]), .CK(i_clk), .RN(n467), .Q(
        inst_r[23]), .QN(n906) );
  DFFRX1 \inst_r_reg[22]  ( .D(inst_w[22]), .CK(i_clk), .RN(n467), .Q(
        inst_r[22]), .QN(n905) );
  DFFRX1 \inst_r_reg[21]  ( .D(inst_w[21]), .CK(i_clk), .RN(n467), .Q(
        inst_r[21]), .QN(n904) );
  DFFRX1 \inst_r_reg[20]  ( .D(inst_w[20]), .CK(i_clk), .RN(n467), .Q(
        inst_r[20]), .QN(n1384) );
  DFFRX1 \inst_r_reg[19]  ( .D(inst_w[19]), .CK(i_clk), .RN(n468), .Q(
        inst_r[19]), .QN(n1385) );
  DFFRX1 \inst_r_reg[18]  ( .D(inst_w[18]), .CK(i_clk), .RN(n468), .Q(
        inst_r[18]), .QN(n1386) );
  DFFRX1 \inst_r_reg[17]  ( .D(inst_w[17]), .CK(i_clk), .RN(n468), .Q(
        inst_r[17]), .QN(n1387) );
  DFFRX1 \inst_r_reg[16]  ( .D(inst_w[16]), .CK(i_clk), .RN(n468), .Q(
        inst_r[16]), .QN(n1388) );
  DFFRX1 ALUSrc_idex_r_reg ( .D(ALUSrc_idex_w), .CK(i_clk), .RN(n469), .Q(n44), 
        .QN(n1389) );
  DFFRX1 \ALUresult2_r_reg[3]  ( .D(n1224), .CK(i_clk), .RN(n462), .QN(n1071)
         );
  DFFRX1 \ALUresult2_r_reg[4]  ( .D(n1222), .CK(i_clk), .RN(n462), .QN(n1069)
         );
  DFFRX1 \ALUresult2_r_reg[5]  ( .D(n1220), .CK(i_clk), .RN(n462), .QN(n1067)
         );
  DFFRX1 \ALUresult2_r_reg[6]  ( .D(n1218), .CK(i_clk), .RN(n462), .QN(n1065)
         );
  DFFRX1 \ALUresult2_r_reg[7]  ( .D(n1216), .CK(i_clk), .RN(n462), .QN(n1063)
         );
  DFFRX1 \ALUresult2_r_reg[8]  ( .D(n1214), .CK(i_clk), .RN(n462), .QN(n1061)
         );
  DFFRX1 \ALUresult2_r_reg[9]  ( .D(n1212), .CK(i_clk), .RN(n462), .QN(n1059)
         );
  DFFRX1 \ALUresult2_r_reg[10]  ( .D(n1210), .CK(i_clk), .RN(n462), .QN(n1057)
         );
  DFFRX1 LO_idex_r_reg ( .D(LO_idex_w), .CK(i_clk), .RN(n466), .QN(n832) );
  DFFRX1 \RegRs_idex_r_reg[4]  ( .D(RegRs_idex_w[4]), .CK(i_clk), .RN(n467), 
        .Q(RegRs_idex_r[4]), .QN(n902) );
  DFFRX1 \RegRs_idex_r_reg[3]  ( .D(RegRs_idex_w[3]), .CK(i_clk), .RN(n467), 
        .Q(RegRs_idex_r[3]), .QN(n901) );
  DFFRX1 \ALUresult2_r_reg[31]  ( .D(n1247), .CK(i_clk), .RN(n465), .QN(n1102)
         );
  DFFRX1 \ALUresult2_r_reg[0]  ( .D(n1245), .CK(i_clk), .RN(n466), .QN(n1100)
         );
  DFFRX1 \ALUresult2_r_reg[1]  ( .D(n1228), .CK(i_clk), .RN(n460), .QN(n1075)
         );
  DFFRX1 \ALUresult2_r_reg[2]  ( .D(n1226), .CK(i_clk), .RN(n460), .QN(n1073)
         );
  DFFRX1 \RegRs_idex_r_reg[2]  ( .D(RegRs_idex_w[2]), .CK(i_clk), .RN(n467), 
        .Q(RegRs_idex_r[2]), .QN(n900) );
  DFFRX1 \RegRs_idex_r_reg[1]  ( .D(RegRs_idex_w[1]), .CK(i_clk), .RN(n467), 
        .Q(RegRs_idex_r[1]), .QN(n899) );
  DFFRX1 \RegRs_idex_r_reg[0]  ( .D(RegRs_idex_w[0]), .CK(i_clk), .RN(n467), 
        .Q(RegRs_idex_r[0]), .QN(n898) );
  DFFRX1 \RegRd_exmem_r_reg[0]  ( .D(n1239), .CK(i_clk), .RN(n466), .Q(
        RegRd_exmem_r[0]), .QN(n1091) );
  DFFRX1 \RegRd_exmem_r_reg[2]  ( .D(n1233), .CK(i_clk), .RN(n460), .Q(
        RegRd_exmem_r[2]), .QN(n1082) );
  DFFRX1 \RegRd_exmem_r_reg[1]  ( .D(n1231), .CK(i_clk), .RN(n460), .Q(
        RegRd_exmem_r[1]), .QN(n1079) );
  DFFRX1 RegWrite_exmem_r_reg ( .D(n1241), .CK(i_clk), .RN(n466), .Q(
        RegWrite_exmem_r), .QN(n1094) );
  DFFRX1 \inst_r_reg[26]  ( .D(inst_w[26]), .CK(i_clk), .RN(n467), .Q(
        inst_r[26]), .QN(n909) );
  DFFRX1 \inst_r_reg[27]  ( .D(inst_w[27]), .CK(i_clk), .RN(n467), .Q(
        inst_r[27]), .QN(n910) );
  DFFRX1 \inst_r_reg[29]  ( .D(inst_w[29]), .CK(i_clk), .RN(n467), .Q(
        inst_r[29]), .QN(n912) );
  DFFRX1 \inst_r_reg[3]  ( .D(inst_w[3]), .CK(i_clk), .RN(n467), .Q(inst_r_3), 
        .QN(n950) );
  DFFRX1 \inst_r_reg[1]  ( .D(inst_w[1]), .CK(i_clk), .RN(n468), .Q(inst_r_1), 
        .QN(n948) );
  DFFRX1 HI_idex_r_reg ( .D(HI_idex_w), .CK(i_clk), .RN(n469), .QN(n799) );
  DFFRX1 Shift_idex_r_reg ( .D(Shift_idex_w), .CK(i_clk), .RN(n466), .Q(n43), 
        .QN(n903) );
  DFFRX1 \ALUresult_r_reg[1]  ( .D(n1229), .CK(i_clk), .RN(n460), .QN(n1428)
         );
  DFFRX1 \ALUresult_r_reg[0]  ( .D(n1246), .CK(i_clk), .RN(n466), .QN(n1429)
         );
  DFFRX1 RegWrite_memwb_r_reg ( .D(n1240), .CK(i_clk), .RN(n466), .Q(
        RegWrite_memwb_r), .QN(n1092) );
  DFFRX1 MemtoReg_memwb_r_reg ( .D(n1249), .CK(i_clk), .RN(n465), .QN(n1105)
         );
  DFFRX1 \RegRd_exmem_r_reg[3]  ( .D(n1235), .CK(i_clk), .RN(n460), .Q(
        RegRd_exmem_r[3]), .QN(n1085) );
  DFFRX1 \RegRd_exmem_r_reg[4]  ( .D(n1237), .CK(i_clk), .RN(n460), .Q(
        RegRd_exmem_r[4]), .QN(n1087) );
  DFFRX1 \RegRt_idex_r_reg[2]  ( .D(RegRt_idex_w[2]), .CK(i_clk), .RN(n468), 
        .Q(RegRt_idex_r[2]), .QN(n1392) );
  DFFRX1 \RegRt_idex_r_reg[0]  ( .D(RegRt_idex_w[0]), .CK(i_clk), .RN(n468), 
        .Q(RegRt_idex_r[0]), .QN(n1394) );
  DFFRX1 \RegRt_idex_r_reg[1]  ( .D(RegRt_idex_w[1]), .CK(i_clk), .RN(n468), 
        .Q(RegRt_idex_r[1]), .QN(n1393) );
  DFFRX1 \RegRt_idex_r_reg[4]  ( .D(RegRt_idex_w[4]), .CK(i_clk), .RN(n467), 
        .Q(RegRt_idex_r[4]), .QN(n1390) );
  DFFRX1 \RegRt_idex_r_reg[3]  ( .D(RegRt_idex_w[3]), .CK(i_clk), .RN(n468), 
        .Q(RegRt_idex_r[3]), .QN(n1391) );
  DFFRX1 \readreg2_2_r_reg[0]  ( .D(n1138), .CK(i_clk), .RN(n469), .Q(n1716), 
        .QN(n954) );
  DFFRX1 \readreg2_2_r_reg[30]  ( .D(n1139), .CK(i_clk), .RN(n468), .Q(n1686), 
        .QN(n956) );
  DFFRX1 \readreg2_2_r_reg[31]  ( .D(n1140), .CK(i_clk), .RN(n474), .Q(n1685), 
        .QN(n958) );
  DFFRX1 \readreg2_2_r_reg[29]  ( .D(n1141), .CK(i_clk), .RN(n474), .Q(n1687), 
        .QN(n960) );
  DFFRX1 \readreg2_2_r_reg[28]  ( .D(n1142), .CK(i_clk), .RN(n474), .Q(n1688), 
        .QN(n962) );
  DFFRX1 \readreg2_2_r_reg[27]  ( .D(n1143), .CK(i_clk), .RN(n474), .Q(n1689), 
        .QN(n964) );
  DFFRX1 \readreg2_2_r_reg[26]  ( .D(n1144), .CK(i_clk), .RN(n474), .Q(n1690), 
        .QN(n966) );
  DFFRX1 \readreg2_2_r_reg[25]  ( .D(n1145), .CK(i_clk), .RN(n474), .Q(n1691), 
        .QN(n968) );
  DFFRX1 \readreg2_2_r_reg[24]  ( .D(n1146), .CK(i_clk), .RN(n474), .Q(n1692), 
        .QN(n970) );
  DFFRX1 \readreg2_2_r_reg[23]  ( .D(n1147), .CK(i_clk), .RN(n474), .Q(n1693), 
        .QN(n972) );
  DFFRX1 \readreg2_2_r_reg[22]  ( .D(n1148), .CK(i_clk), .RN(n474), .Q(n1694), 
        .QN(n974) );
  DFFRX1 \readreg2_2_r_reg[21]  ( .D(n1149), .CK(i_clk), .RN(n474), .Q(n1695), 
        .QN(n976) );
  DFFRX1 \readreg2_2_r_reg[20]  ( .D(n1150), .CK(i_clk), .RN(n474), .Q(n1696), 
        .QN(n978) );
  DFFRX1 \readreg2_2_r_reg[19]  ( .D(n1151), .CK(i_clk), .RN(n474), .Q(n1697), 
        .QN(n980) );
  DFFRX1 \readreg2_2_r_reg[18]  ( .D(n1152), .CK(i_clk), .RN(n474), .Q(n1698), 
        .QN(n982) );
  DFFRX1 \readreg2_2_r_reg[17]  ( .D(n1153), .CK(i_clk), .RN(n474), .Q(n1699), 
        .QN(n984) );
  DFFRX1 \readreg2_2_r_reg[16]  ( .D(n1154), .CK(i_clk), .RN(n474), .Q(n1700), 
        .QN(n986) );
  DFFRX1 \readreg2_2_r_reg[15]  ( .D(n1155), .CK(i_clk), .RN(n473), .Q(n1701), 
        .QN(n988) );
  DFFRX1 \readreg2_2_r_reg[14]  ( .D(n1156), .CK(i_clk), .RN(n473), .Q(n1702), 
        .QN(n990) );
  DFFRX1 \readreg2_2_r_reg[13]  ( .D(n1157), .CK(i_clk), .RN(n473), .Q(n1703), 
        .QN(n992) );
  DFFRX1 \readreg2_2_r_reg[12]  ( .D(n1158), .CK(i_clk), .RN(n473), .Q(n1704), 
        .QN(n994) );
  DFFRX1 \readreg2_2_r_reg[11]  ( .D(n1159), .CK(i_clk), .RN(n473), .Q(n1705), 
        .QN(n996) );
  DFFRX1 \readreg2_2_r_reg[10]  ( .D(n1160), .CK(i_clk), .RN(n473), .Q(n1706), 
        .QN(n998) );
  DFFRX1 \readreg2_2_r_reg[9]  ( .D(n1161), .CK(i_clk), .RN(n473), .Q(n1707), 
        .QN(n1000) );
  DFFRX1 \readreg2_2_r_reg[8]  ( .D(n1162), .CK(i_clk), .RN(n473), .Q(n1708), 
        .QN(n1002) );
  DFFRX1 \readreg2_2_r_reg[7]  ( .D(n1163), .CK(i_clk), .RN(n473), .Q(n1709), 
        .QN(n1004) );
  DFFRX1 \readreg2_2_r_reg[6]  ( .D(n1164), .CK(i_clk), .RN(n473), .Q(n1710), 
        .QN(n1006) );
  DFFRX1 \readreg2_2_r_reg[5]  ( .D(n1165), .CK(i_clk), .RN(n473), .Q(n1711), 
        .QN(n1008) );
  DFFRX1 \readreg2_2_r_reg[4]  ( .D(n1166), .CK(i_clk), .RN(n473), .Q(n1712), 
        .QN(n1010) );
  DFFRX1 \readreg2_2_r_reg[3]  ( .D(n1167), .CK(i_clk), .RN(n473), .Q(n1713), 
        .QN(n1012) );
  DFFRX1 \readreg2_2_r_reg[2]  ( .D(n1168), .CK(i_clk), .RN(n473), .Q(n1714), 
        .QN(n1014) );
  DFFRX1 \readreg2_2_r_reg[1]  ( .D(n1169), .CK(i_clk), .RN(n473), .Q(n1715), 
        .QN(n1016) );
  DFFRX1 \ALUresult_r_reg[6]  ( .D(n1219), .CK(i_clk), .RN(n462), .Q(n1684), 
        .QN(n1423) );
  DFFRX1 \RegRd_memwb_r_reg[2]  ( .D(n1232), .CK(i_clk), .RN(n460), .Q(
        RegRd_memwb_r[2]), .QN(n1080) );
  DFFRX1 \RegRd_memwb_r_reg[1]  ( .D(n1230), .CK(i_clk), .RN(n460), .Q(
        RegRd_memwb_r[1]), .QN(n1077) );
  DFFRX1 \RegRd_memwb_r_reg[3]  ( .D(n1234), .CK(i_clk), .RN(n460), .Q(
        RegRd_memwb_r[3]), .QN(n1083) );
  DFFRX1 \inst_r_reg[31]  ( .D(inst_w[31]), .CK(i_clk), .RN(n467), .QN(n914)
         );
  DFFRX1 \readdata_r_reg[30]  ( .D(n1280), .CK(i_clk), .RN(n466), .Q(n1136) );
  DFFRX1 \readdata_r_reg[29]  ( .D(n1279), .CK(i_clk), .RN(n465), .Q(n1135) );
  DFFRX1 \readdata_r_reg[28]  ( .D(n1278), .CK(i_clk), .RN(n465), .Q(n1134) );
  DFFRX1 \readdata_r_reg[27]  ( .D(n1277), .CK(i_clk), .RN(n465), .Q(n1133) );
  DFFRX1 \readdata_r_reg[26]  ( .D(n1276), .CK(i_clk), .RN(n465), .Q(n1132) );
  DFFRX1 \readdata_r_reg[25]  ( .D(n1275), .CK(i_clk), .RN(n465), .Q(n1131) );
  DFFRX1 \readdata_r_reg[24]  ( .D(n1274), .CK(i_clk), .RN(n465), .Q(n1130) );
  DFFRX1 \readdata_r_reg[23]  ( .D(n1273), .CK(i_clk), .RN(n465), .Q(n1129) );
  DFFRX1 \readdata_r_reg[22]  ( .D(n1272), .CK(i_clk), .RN(n465), .Q(n1128) );
  DFFRX1 \readdata_r_reg[21]  ( .D(n1271), .CK(i_clk), .RN(n465), .Q(n1127) );
  DFFRX1 \readdata_r_reg[20]  ( .D(n1270), .CK(i_clk), .RN(n465), .Q(n1126) );
  DFFRX1 \readdata_r_reg[19]  ( .D(n1269), .CK(i_clk), .RN(n465), .Q(n1125) );
  DFFRX1 \readdata_r_reg[18]  ( .D(n1268), .CK(i_clk), .RN(n465), .Q(n1124) );
  DFFRX1 \readdata_r_reg[17]  ( .D(n1267), .CK(i_clk), .RN(n465), .Q(n1123) );
  DFFRX1 \readdata_r_reg[16]  ( .D(n1266), .CK(i_clk), .RN(n465), .Q(n1122) );
  DFFRX1 \readdata_r_reg[6]  ( .D(n1256), .CK(i_clk), .RN(n465), .Q(n1112) );
  DFFRX1 \readdata_r_reg[31]  ( .D(n1281), .CK(i_clk), .RN(n468), .Q(n1137) );
  DFFRX1 \readdata_r_reg[15]  ( .D(n1265), .CK(i_clk), .RN(n465), .Q(n1121) );
  DFFRX1 \readdata_r_reg[14]  ( .D(n1264), .CK(i_clk), .RN(n465), .Q(n1120) );
  DFFRX1 \readdata_r_reg[13]  ( .D(n1263), .CK(i_clk), .RN(n465), .Q(n1119) );
  DFFRX1 \readdata_r_reg[12]  ( .D(n1262), .CK(i_clk), .RN(n465), .Q(n1118) );
  DFFRX1 \readdata_r_reg[11]  ( .D(n1261), .CK(i_clk), .RN(n465), .Q(n1117) );
  DFFRX1 \readdata_r_reg[10]  ( .D(n1260), .CK(i_clk), .RN(n465), .Q(n1116) );
  DFFRX1 \readdata_r_reg[9]  ( .D(n1259), .CK(i_clk), .RN(n465), .Q(n1115) );
  DFFRX1 \readdata_r_reg[8]  ( .D(n1258), .CK(i_clk), .RN(n465), .Q(n1114) );
  DFFRX1 \readdata_r_reg[7]  ( .D(n1257), .CK(i_clk), .RN(n465), .Q(n1113) );
  DFFRX1 \readdata_r_reg[5]  ( .D(n1255), .CK(i_clk), .RN(n465), .Q(n1111) );
  DFFRX1 \readdata_r_reg[4]  ( .D(n1254), .CK(i_clk), .RN(n465), .Q(n1110) );
  DFFRX1 \readdata_r_reg[3]  ( .D(n1253), .CK(i_clk), .RN(n465), .Q(n1109) );
  DFFRX1 \readdata_r_reg[2]  ( .D(n1252), .CK(i_clk), .RN(n465), .Q(n1108) );
  DFFRX1 \readdata_r_reg[1]  ( .D(n1251), .CK(i_clk), .RN(n465), .Q(n1107) );
  DFFRX1 \readdata_r_reg[0]  ( .D(n1250), .CK(i_clk), .RN(n465), .Q(n1106) );
  DFFRX1 \shamt_idex_r_reg[4]  ( .D(shamt_idex_w[4]), .CK(i_clk), .RN(n460), 
        .Q(shamt_idex_r[4]) );
  DFFRX1 \shamt_idex_r_reg[3]  ( .D(shamt_idex_w[3]), .CK(i_clk), .RN(n466), 
        .Q(shamt_idex_r[3]) );
  DFFRX1 \shamt_idex_r_reg[0]  ( .D(shamt_idex_w[0]), .CK(i_clk), .RN(n466), 
        .Q(shamt_idex_r[0]) );
  DFFRX1 \shamt_idex_r_reg[2]  ( .D(shamt_idex_w[2]), .CK(i_clk), .RN(n466), 
        .Q(shamt_idex_r[2]) );
  DFFRX1 \shamt_idex_r_reg[1]  ( .D(shamt_idex_w[1]), .CK(i_clk), .RN(n466), 
        .Q(shamt_idex_r[1]) );
  DFFRX1 \sign_ext_r_reg[8]  ( .D(sign_ext_w[8]), .CK(i_clk), .RN(n466), .QN(
        n1542) );
  DFFRX1 \readreg1_r_reg[16]  ( .D(readreg1_w[16]), .CK(i_clk), .RN(n468), 
        .QN(n1628) );
  DFFRX1 \readreg1_r_reg[15]  ( .D(readreg1_w[15]), .CK(i_clk), .RN(n470), 
        .QN(n1627) );
  DFFRX1 \readreg1_r_reg[14]  ( .D(readreg1_w[14]), .CK(i_clk), .RN(n475), 
        .QN(n1626) );
  DFFRX1 \readreg1_r_reg[13]  ( .D(readreg1_w[13]), .CK(i_clk), .RN(n475), 
        .QN(n1625) );
  DFFRX1 \readreg1_r_reg[12]  ( .D(readreg1_w[12]), .CK(i_clk), .RN(n475), 
        .QN(n1624) );
  DFFRX1 \readreg1_r_reg[11]  ( .D(readreg1_w[11]), .CK(i_clk), .RN(n475), 
        .QN(n1623) );
  DFFRX1 \readreg1_r_reg[10]  ( .D(readreg1_w[10]), .CK(i_clk), .RN(n475), 
        .QN(n1622) );
  DFFRX1 \readreg1_r_reg[0]  ( .D(readreg1_w[0]), .CK(i_clk), .RN(n474), .QN(
        n1612) );
  DFFRX1 \sign_ext_r_reg[11]  ( .D(sign_ext_w[11]), .CK(i_clk), .RN(n466), 
        .QN(n1537) );
  DFFRX1 \sign_ext_r_reg[10]  ( .D(sign_ext_w[10]), .CK(i_clk), .RN(n460), 
        .QN(n1577) );
  DFFRX1 \sign_ext_r_reg[9]  ( .D(sign_ext_w[9]), .CK(i_clk), .RN(n466), .QN(
        n1540) );
  DFFRX1 \sign_ext_r_reg[5]  ( .D(sign_ext_w[5]), .CK(i_clk), .RN(n467), .QN(
        n1547) );
  DFFRX1 \sign_ext_r_reg[4]  ( .D(sign_ext_w[4]), .CK(i_clk), .RN(n467), .QN(
        n1548) );
  DFFRX1 \sign_ext_r_reg[3]  ( .D(sign_ext_w[3]), .CK(i_clk), .RN(n467), .QN(
        n1549) );
  DFFRX1 \sign_ext_r_reg[2]  ( .D(sign_ext_w[2]), .CK(i_clk), .RN(n467), .QN(
        n1551) );
  DFFRX1 \sign_ext_r_reg[1]  ( .D(sign_ext_w[1]), .CK(i_clk), .RN(n468), .QN(
        n1552) );
  DFFRX1 \sign_ext_r_reg[0]  ( .D(sign_ext_w[0]), .CK(i_clk), .RN(n460), .QN(
        n1578) );
  DFFRX1 \readreg2_r_reg[31]  ( .D(readreg2_w[31]), .CK(i_clk), .RN(n474), 
        .QN(n1611) );
  DFFRX1 \readreg2_r_reg[30]  ( .D(readreg2_w[30]), .CK(i_clk), .RN(n474), 
        .QN(n1610) );
  DFFRX1 \readreg2_r_reg[29]  ( .D(readreg2_w[29]), .CK(i_clk), .RN(n474), 
        .QN(n1609) );
  DFFRX1 \readreg2_r_reg[28]  ( .D(readreg2_w[28]), .CK(i_clk), .RN(n474), 
        .QN(n1608) );
  DFFRX1 \readreg2_r_reg[27]  ( .D(readreg2_w[27]), .CK(i_clk), .RN(n474), 
        .QN(n1607) );
  DFFRX1 \readreg2_r_reg[26]  ( .D(readreg2_w[26]), .CK(i_clk), .RN(n474), 
        .QN(n1606) );
  DFFRX1 \readreg2_r_reg[25]  ( .D(readreg2_w[25]), .CK(i_clk), .RN(n474), 
        .QN(n1605) );
  DFFRX1 \readreg2_r_reg[24]  ( .D(readreg2_w[24]), .CK(i_clk), .RN(n474), 
        .QN(n1604) );
  DFFRX1 \readreg2_r_reg[23]  ( .D(readreg2_w[23]), .CK(i_clk), .RN(n474), 
        .QN(n1603) );
  DFFRX1 \readreg2_r_reg[22]  ( .D(readreg2_w[22]), .CK(i_clk), .RN(n474), 
        .QN(n1602) );
  DFFRX1 \readreg2_r_reg[21]  ( .D(readreg2_w[21]), .CK(i_clk), .RN(n474), 
        .QN(n1601) );
  DFFRX1 \readreg2_r_reg[20]  ( .D(readreg2_w[20]), .CK(i_clk), .RN(n474), 
        .QN(n1600) );
  DFFRX1 \readreg2_r_reg[19]  ( .D(readreg2_w[19]), .CK(i_clk), .RN(n474), 
        .QN(n1599) );
  DFFRX1 \readreg2_r_reg[18]  ( .D(readreg2_w[18]), .CK(i_clk), .RN(n474), 
        .QN(n1598) );
  DFFRX1 \readreg2_r_reg[16]  ( .D(readreg2_w[16]), .CK(i_clk), .RN(n473), 
        .QN(n1596) );
  DFFRX1 \readreg2_r_reg[13]  ( .D(readreg2_w[13]), .CK(i_clk), .RN(n473), 
        .QN(n1593) );
  DFFRX1 \readreg2_r_reg[10]  ( .D(readreg2_w[10]), .CK(i_clk), .RN(n473), 
        .QN(n1590) );
  DFFRX1 \readreg2_r_reg[9]  ( .D(readreg2_w[9]), .CK(i_clk), .RN(n473), .QN(
        n1589) );
  DFFRX1 \readreg2_r_reg[8]  ( .D(readreg2_w[8]), .CK(i_clk), .RN(n473), .QN(
        n1588) );
  DFFRX1 \readreg2_r_reg[7]  ( .D(readreg2_w[7]), .CK(i_clk), .RN(n473), .QN(
        n1587) );
  DFFRX1 \readreg2_r_reg[6]  ( .D(readreg2_w[6]), .CK(i_clk), .RN(n473), .QN(
        n1586) );
  DFFRX1 \readreg2_r_reg[5]  ( .D(readreg2_w[5]), .CK(i_clk), .RN(n473), .QN(
        n1585) );
  DFFRX1 \readreg2_r_reg[4]  ( .D(readreg2_w[4]), .CK(i_clk), .RN(n473), .QN(
        n1584) );
  DFFRX1 \readreg2_r_reg[3]  ( .D(readreg2_w[3]), .CK(i_clk), .RN(n473), .QN(
        n1583) );
  DFFRX1 \readreg2_r_reg[2]  ( .D(readreg2_w[2]), .CK(i_clk), .RN(n473), .QN(
        n1582) );
  DFFRX1 \readreg2_r_reg[1]  ( .D(readreg2_w[1]), .CK(i_clk), .RN(n473), .QN(
        n1581) );
  DFFRX1 \readreg2_r_reg[0]  ( .D(readreg2_w[0]), .CK(i_clk), .RN(n473), .QN(
        n1580) );
  DFFRX1 \readreg1_r_reg[31]  ( .D(readreg1_w[31]), .CK(i_clk), .RN(n468), 
        .QN(n1643) );
  DFFRX1 \readreg1_r_reg[30]  ( .D(readreg1_w[30]), .CK(i_clk), .RN(n468), 
        .QN(n1642) );
  DFFRX1 \readreg1_r_reg[29]  ( .D(readreg1_w[29]), .CK(i_clk), .RN(n468), 
        .QN(n1641) );
  DFFRX1 \readreg1_r_reg[28]  ( .D(readreg1_w[28]), .CK(i_clk), .RN(n468), 
        .QN(n1640) );
  DFFRX1 \readreg1_r_reg[27]  ( .D(readreg1_w[27]), .CK(i_clk), .RN(n468), 
        .QN(n1639) );
  DFFRX1 \readreg1_r_reg[26]  ( .D(readreg1_w[26]), .CK(i_clk), .RN(n468), 
        .QN(n1638) );
  DFFRX1 \readreg1_r_reg[25]  ( .D(readreg1_w[25]), .CK(i_clk), .RN(n468), 
        .QN(n1637) );
  DFFRX1 \readreg1_r_reg[24]  ( .D(readreg1_w[24]), .CK(i_clk), .RN(n468), 
        .QN(n1636) );
  DFFRX1 \readreg1_r_reg[23]  ( .D(readreg1_w[23]), .CK(i_clk), .RN(n468), 
        .QN(n1635) );
  DFFRX1 \readreg1_r_reg[22]  ( .D(readreg1_w[22]), .CK(i_clk), .RN(n468), 
        .QN(n1634) );
  DFFRX1 \readreg1_r_reg[21]  ( .D(readreg1_w[21]), .CK(i_clk), .RN(n468), 
        .QN(n1633) );
  DFFRX1 \readreg1_r_reg[20]  ( .D(readreg1_w[20]), .CK(i_clk), .RN(n468), 
        .QN(n1632) );
  DFFRX1 \readreg1_r_reg[19]  ( .D(readreg1_w[19]), .CK(i_clk), .RN(n468), 
        .QN(n1631) );
  DFFRX1 \readreg1_r_reg[18]  ( .D(readreg1_w[18]), .CK(i_clk), .RN(n468), 
        .QN(n1630) );
  DFFRX1 \readreg1_r_reg[17]  ( .D(readreg1_w[17]), .CK(i_clk), .RN(n468), 
        .QN(n1629) );
  DFFRX1 \readreg1_r_reg[9]  ( .D(readreg1_w[9]), .CK(i_clk), .RN(n475), .QN(
        n1621) );
  DFFRX1 \readreg1_r_reg[8]  ( .D(readreg1_w[8]), .CK(i_clk), .RN(n475), .QN(
        n1620) );
  DFFRX1 \readreg1_r_reg[7]  ( .D(readreg1_w[7]), .CK(i_clk), .RN(n475), .QN(
        n1619) );
  DFFRX1 \readreg1_r_reg[6]  ( .D(readreg1_w[6]), .CK(i_clk), .RN(n475), .QN(
        n1618) );
  DFFRX1 \readreg1_r_reg[5]  ( .D(readreg1_w[5]), .CK(i_clk), .RN(n475), .QN(
        n1617) );
  DFFRX1 \readreg1_r_reg[4]  ( .D(readreg1_w[4]), .CK(i_clk), .RN(n474), .QN(
        n1616) );
  DFFRX1 \readreg1_r_reg[3]  ( .D(readreg1_w[3]), .CK(i_clk), .RN(n474), .QN(
        n1615) );
  DFFRX1 \readreg1_r_reg[2]  ( .D(readreg1_w[2]), .CK(i_clk), .RN(n474), .QN(
        n1614) );
  DFFRX1 \readreg1_r_reg[1]  ( .D(readreg1_w[1]), .CK(i_clk), .RN(n474), .QN(
        n1613) );
  DFFRX1 \readreg2_r_reg[17]  ( .D(readreg2_w[17]), .CK(i_clk), .RN(n474), 
        .QN(n1597) );
  DFFRX1 \readreg2_r_reg[15]  ( .D(readreg2_w[15]), .CK(i_clk), .RN(n473), 
        .QN(n1595) );
  DFFRX1 \readreg2_r_reg[14]  ( .D(readreg2_w[14]), .CK(i_clk), .RN(n473), 
        .QN(n1594) );
  DFFRX1 \readreg2_r_reg[12]  ( .D(readreg2_w[12]), .CK(i_clk), .RN(n473), 
        .QN(n1592) );
  DFFRX1 \readreg2_r_reg[11]  ( .D(readreg2_w[11]), .CK(i_clk), .RN(n473), 
        .QN(n1591) );
  DFFRX1 \sign_ext_r_reg[14]  ( .D(sign_ext_w[14]), .CK(i_clk), .RN(n460), 
        .QN(n1571) );
  DFFRX1 \sign_ext_r_reg[13]  ( .D(sign_ext_w[13]), .CK(i_clk), .RN(n460), 
        .QN(n1573) );
  DFFRX1 \sign_ext_r_reg[12]  ( .D(sign_ext_w[12]), .CK(i_clk), .RN(n460), 
        .QN(n1575) );
  DFFRX1 \sign_ext_r_reg[7]  ( .D(sign_ext_w[7]), .CK(i_clk), .RN(n466), .QN(
        n1544) );
  DFFRX1 \sign_ext_r_reg[6]  ( .D(sign_ext_w[6]), .CK(i_clk), .RN(n466), .QN(
        n1546) );
  DFFRX1 \ALUOp_idex_r_reg[0]  ( .D(ALUOp_idex_w[0]), .CK(i_clk), .RN(n470), 
        .Q(ALUOp_idex_r[0]) );
  DFFRX1 \ALUOp_idex_r_reg[1]  ( .D(ALUOp_idex_w[1]), .CK(i_clk), .RN(n470), 
        .Q(ALUOp_idex_r[1]) );
  DFFRX1 \sign_ext_r_reg[31]  ( .D(sign_ext_w[31]), .CK(i_clk), .RN(n468), 
        .QN(n1553) );
  DFFRX1 \sign_ext_r_reg[30]  ( .D(sign_ext_w[30]), .CK(i_clk), .RN(n468), 
        .QN(n1554) );
  DFFRX1 \sign_ext_r_reg[29]  ( .D(sign_ext_w[29]), .CK(i_clk), .RN(n468), 
        .QN(n1555) );
  DFFRX1 \sign_ext_r_reg[28]  ( .D(sign_ext_w[28]), .CK(i_clk), .RN(n462), 
        .QN(n1556) );
  DFFRX1 \sign_ext_r_reg[27]  ( .D(sign_ext_w[27]), .CK(i_clk), .RN(n458), 
        .QN(n1557) );
  DFFRX1 \sign_ext_r_reg[26]  ( .D(sign_ext_w[26]), .CK(i_clk), .RN(n458), 
        .QN(n1558) );
  DFFRX1 \sign_ext_r_reg[25]  ( .D(sign_ext_w[25]), .CK(i_clk), .RN(n458), 
        .QN(n1559) );
  DFFRX1 \sign_ext_r_reg[24]  ( .D(sign_ext_w[24]), .CK(i_clk), .RN(n458), 
        .QN(n1560) );
  DFFRX1 \sign_ext_r_reg[23]  ( .D(sign_ext_w[23]), .CK(i_clk), .RN(n458), 
        .QN(n1561) );
  DFFRX1 \sign_ext_r_reg[22]  ( .D(sign_ext_w[22]), .CK(i_clk), .RN(n458), 
        .QN(n1562) );
  DFFRX1 \sign_ext_r_reg[21]  ( .D(sign_ext_w[21]), .CK(i_clk), .RN(n458), 
        .QN(n1563) );
  DFFRX1 \sign_ext_r_reg[20]  ( .D(sign_ext_w[20]), .CK(i_clk), .RN(n458), 
        .QN(n1564) );
  DFFRX1 \sign_ext_r_reg[19]  ( .D(sign_ext_w[19]), .CK(i_clk), .RN(n458), 
        .QN(n1565) );
  DFFRX1 \sign_ext_r_reg[18]  ( .D(sign_ext_w[18]), .CK(i_clk), .RN(n458), 
        .QN(n1566) );
  DFFRX1 \sign_ext_r_reg[17]  ( .D(sign_ext_w[17]), .CK(i_clk), .RN(n458), 
        .QN(n1567) );
  DFFRX1 \sign_ext_r_reg[16]  ( .D(sign_ext_w[16]), .CK(i_clk), .RN(n458), 
        .QN(n1568) );
  DFFRX1 \sign_ext_r_reg[15]  ( .D(sign_ext_w[15]), .CK(i_clk), .RN(n458), 
        .QN(n1569) );
  DFFRX1 \inst_r_reg[8]  ( .D(inst_w[8]), .CK(i_clk), .RN(n466), .Q(
        sign_ext[8]), .QN(n1541) );
  DFFRX1 \inst_r_reg[7]  ( .D(inst_w[7]), .CK(i_clk), .RN(n466), .Q(
        sign_ext[7]), .QN(n1543) );
  DFFRX1 \inst_r_reg[6]  ( .D(inst_w[6]), .CK(i_clk), .RN(n466), .Q(
        sign_ext[6]), .QN(n1545) );
  DFFRX1 \inst_r_reg[9]  ( .D(inst_w[9]), .CK(i_clk), .RN(n466), .Q(
        sign_ext[9]), .QN(n1539) );
  DFFRX1 take_r_reg ( .D(take_w), .CK(i_clk), .RN(n466), .Q(take_r), .QN(n1538) );
  DFFRX1 \inst_r_reg[15]  ( .D(inst_w[15]), .CK(i_clk), .RN(n468), .Q(
        sign_ext_31), .QN(n45) );
  DFFRX1 \inst_r_reg[14]  ( .D(inst_w[14]), .CK(i_clk), .RN(n460), .Q(
        sign_ext[14]), .QN(n1570) );
  DFFRX1 \inst_r_reg[13]  ( .D(inst_w[13]), .CK(i_clk), .RN(n460), .Q(
        sign_ext[13]), .QN(n1572) );
  DFFRX1 \inst_r_reg[12]  ( .D(inst_w[12]), .CK(i_clk), .RN(n460), .Q(
        sign_ext[12]), .QN(n1574) );
  DFFRX1 \inst_r_reg[11]  ( .D(inst_w[11]), .CK(i_clk), .RN(n466), .Q(
        sign_ext[11]), .QN(n1536) );
  DFFRX1 \inst_r_reg[10]  ( .D(inst_w[10]), .CK(i_clk), .RN(n460), .Q(
        sign_ext[10]), .QN(n1576) );
  DFFRX1 \PC_r_reg[0]  ( .D(PC_w[0]), .CK(i_clk), .RN(n460), .Q(PC_r[0]), .QN(
        n1579) );
  DFFRX1 \PC_r_reg[8]  ( .D(PC_w[8]), .CK(i_clk), .RN(n469), .Q(ICACHE_addr[6]) );
  DFFRX1 \PC_r_reg[1]  ( .D(PC_w[1]), .CK(i_clk), .RN(n468), .Q(PC_r[1]), .QN(
        n644) );
  DFFRX1 \PC_r_reg[7]  ( .D(PC_w[7]), .CK(i_clk), .RN(n469), .Q(ICACHE_addr[5]) );
  DFFRX1 \PC_r_reg[6]  ( .D(PC_w[6]), .CK(i_clk), .RN(n469), .Q(ICACHE_addr[4]) );
  DFFRX1 \PC_r_reg[3]  ( .D(PC_w[3]), .CK(i_clk), .RN(n469), .Q(ICACHE_addr[1]) );
  DFFRX1 \PC_r_reg[14]  ( .D(PC_w[14]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[12]) );
  DFFRX1 \PC_r_reg[11]  ( .D(PC_w[11]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[9]) );
  DFFRX1 \PC_r_reg[13]  ( .D(PC_w[13]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[11]) );
  DFFRX1 \PC_r_reg[12]  ( .D(PC_w[12]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[10]) );
  DFFRX1 \PC_r_reg[10]  ( .D(PC_w[10]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[8]) );
  DFFRX1 \PC_r_reg[9]  ( .D(PC_w[9]), .CK(i_clk), .RN(n469), .Q(ICACHE_addr[7]) );
  DFFRX1 \PC_r_reg[15]  ( .D(PC_w[15]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[13]) );
  DFFRX1 \PC_r_reg[16]  ( .D(PC_w[16]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[14]) );
  DFFRX1 \PC_r_reg[17]  ( .D(PC_w[17]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[15]) );
  DFFRX1 \PC_r_reg[18]  ( .D(PC_w[18]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[16]) );
  DFFRX1 \PC_r_reg[19]  ( .D(PC_w[19]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[17]) );
  DFFRX1 \PC_r_reg[20]  ( .D(PC_w[20]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[18]) );
  DFFRX1 \PC_r_reg[21]  ( .D(PC_w[21]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[19]) );
  DFFRX1 \PC_r_reg[22]  ( .D(PC_w[22]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[20]) );
  DFFRX1 \PC_r_reg[23]  ( .D(PC_w[23]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[21]) );
  DFFRX1 \PC_r_reg[24]  ( .D(PC_w[24]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[22]) );
  DFFRX1 \PC_r_reg[25]  ( .D(PC_w[25]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[23]) );
  DFFRX1 \PC_r_reg[26]  ( .D(PC_w[26]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[24]) );
  DFFRX1 \PC_r_reg[27]  ( .D(PC_w[27]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[25]) );
  DFFRX1 \PC_r_reg[28]  ( .D(PC_w[28]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[26]) );
  DFFRX1 \PC_r_reg[29]  ( .D(PC_w[29]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[27]) );
  DFFRX1 \PC_r_reg[30]  ( .D(PC_w[30]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[28]) );
  DFFRX1 \PC_r_reg[31]  ( .D(PC_w[31]), .CK(i_clk), .RN(n469), .Q(
        ICACHE_addr[29]) );
  DFFRX1 MemWrite_exmem_r_reg ( .D(n1242), .CK(i_clk), .RN(n466), .QN(n1096)
         );
  DFFRX1 \ALUresult_r_reg[4]  ( .D(n1223), .CK(i_clk), .RN(n462), .Q(n184), 
        .QN(n1425) );
  DFFRX1 \ALUresult_r_reg[5]  ( .D(n1221), .CK(i_clk), .RN(n462), .Q(n141), 
        .QN(n1424) );
  DFFRX1 \ALUresult_r_reg[3]  ( .D(n1225), .CK(i_clk), .RN(n462), .Q(n140), 
        .QN(n1426) );
  DFFRX1 \ALUresult_r_reg[2]  ( .D(n1227), .CK(i_clk), .RN(n460), .Q(n183), 
        .QN(n1427) );
  DFFRX1 \ALUresult_r_reg[7]  ( .D(n1217), .CK(i_clk), .RN(n462), .Q(n144), 
        .QN(n1422) );
  DFFRX1 \ALUresult_r_reg[8]  ( .D(n1215), .CK(i_clk), .RN(n462), .Q(n191), 
        .QN(n1421) );
  DFFRX1 \ALUresult_r_reg[9]  ( .D(n1213), .CK(i_clk), .RN(n462), .Q(n135), 
        .QN(n1420) );
  DFFRX1 \ALUresult_r_reg[10]  ( .D(n1211), .CK(i_clk), .RN(n462), .Q(n185), 
        .QN(n1419) );
  DFFRX1 \ALUresult_r_reg[11]  ( .D(n1209), .CK(i_clk), .RN(n464), .Q(n143), 
        .QN(n1418) );
  DFFRX1 \ALUresult_r_reg[12]  ( .D(n1207), .CK(i_clk), .RN(n464), .Q(n139), 
        .QN(n1417) );
  DFFRX1 \ALUresult_r_reg[13]  ( .D(n1205), .CK(i_clk), .RN(n464), .Q(n188), 
        .QN(n1416) );
  DFFRX1 \ALUresult_r_reg[14]  ( .D(n1203), .CK(i_clk), .RN(n464), .Q(n137), 
        .QN(n1415) );
  DFFRX1 \ALUresult_r_reg[15]  ( .D(n1201), .CK(i_clk), .RN(n464), .Q(n147), 
        .QN(n1414) );
  DFFRX1 \ALUresult_r_reg[16]  ( .D(n1199), .CK(i_clk), .RN(n464), .Q(n193), 
        .QN(n1413) );
  DFFRX1 \ALUresult_r_reg[17]  ( .D(n1197), .CK(i_clk), .RN(n464), .Q(n149), 
        .QN(n1412) );
  DFFRX1 \ALUresult_r_reg[18]  ( .D(n1195), .CK(i_clk), .RN(n464), .Q(n195), 
        .QN(n1411) );
  DFFRX1 \ALUresult_r_reg[19]  ( .D(n1193), .CK(i_clk), .RN(n464), .Q(n136), 
        .QN(n1410) );
  DFFRX1 \ALUresult_r_reg[20]  ( .D(n1191), .CK(i_clk), .RN(n473), .Q(n134), 
        .QN(n1409) );
  DFFRX1 \ALUresult_r_reg[21]  ( .D(n1189), .CK(i_clk), .RN(n471), .Q(n142), 
        .QN(n1408) );
  DFFRX1 \ALUresult_r_reg[22]  ( .D(n1187), .CK(i_clk), .RN(n472), .Q(n186), 
        .QN(n1407) );
  DFFRX1 \ALUresult_r_reg[23]  ( .D(n1185), .CK(i_clk), .RN(n472), .Q(n190), 
        .QN(n1406) );
  DFFRX1 \ALUresult_r_reg[24]  ( .D(n1183), .CK(i_clk), .RN(n472), .Q(n187), 
        .QN(n1405) );
  DFFRX1 \ALUresult_r_reg[25]  ( .D(n1181), .CK(i_clk), .RN(n472), .Q(n145), 
        .QN(n1404) );
  DFFRX1 \ALUresult_r_reg[26]  ( .D(n1179), .CK(i_clk), .RN(n472), .Q(n138), 
        .QN(n1403) );
  DFFRX1 \ALUresult_r_reg[27]  ( .D(n1177), .CK(i_clk), .RN(n472), .Q(n148), 
        .QN(n1402) );
  DFFRX1 \ALUresult_r_reg[28]  ( .D(n1175), .CK(i_clk), .RN(n472), .Q(n194), 
        .QN(n1401) );
  DFFRX1 \ALUresult_r_reg[29]  ( .D(n1173), .CK(i_clk), .RN(n472), .Q(n146), 
        .QN(n1400) );
  DFFRX1 \ALUresult_r_reg[30]  ( .D(n1171), .CK(i_clk), .RN(n473), .Q(n192), 
        .QN(n1399) );
  DFFRX1 \ALUresult_r_reg[31]  ( .D(n1248), .CK(i_clk), .RN(n465), .Q(n133), 
        .QN(n1398) );
  DFFRX1 \LO_r_reg[7]  ( .D(n923), .CK(i_clk), .RN(n470), .Q(n1651), .QN(n862)
         );
  DFFRX1 \LO_r_reg[6]  ( .D(n924), .CK(i_clk), .RN(n470), .Q(n1650), .QN(n861)
         );
  DFFRX1 \LO_r_reg[8]  ( .D(n922), .CK(i_clk), .RN(n470), .Q(n1652), .QN(n863)
         );
  DFFRX1 \HI_r_reg[0]  ( .D(n1287), .CK(i_clk), .RN(n471), .Q(n1664), .QN(n800) );
  DFFRX1 \LO_r_reg[1]  ( .D(n941), .CK(i_clk), .RN(n470), .Q(n1645), .QN(n844)
         );
  DFFRX1 \LO_r_reg[0]  ( .D(n963), .CK(i_clk), .RN(n470), .Q(n1644), .QN(n833)
         );
  DFFRX1 \HI_r_reg[8]  ( .D(n967), .CK(i_clk), .RN(n471), .Q(n1672), .QN(n830)
         );
  DFFRX1 \HI_r_reg[7]  ( .D(n969), .CK(i_clk), .RN(n471), .Q(n1671), .QN(n829)
         );
  DFFRX1 \HI_r_reg[6]  ( .D(n971), .CK(i_clk), .RN(n471), .Q(n1670), .QN(n828)
         );
  DFFRX1 \HI_r_reg[5]  ( .D(n973), .CK(i_clk), .RN(n471), .Q(n1669), .QN(n827)
         );
  DFFRX1 \HI_r_reg[4]  ( .D(n975), .CK(i_clk), .RN(n471), .Q(n1668), .QN(n826)
         );
  DFFRX1 \HI_r_reg[3]  ( .D(n977), .CK(i_clk), .RN(n471), .Q(n1667), .QN(n825)
         );
  DFFRX1 \HI_r_reg[2]  ( .D(n983), .CK(i_clk), .RN(n471), .Q(n1666), .QN(n822)
         );
  DFFRX1 \HI_r_reg[1]  ( .D(n1005), .CK(i_clk), .RN(n471), .Q(n1665), .QN(n811) );
  DFFRX1 \LO_r_reg[5]  ( .D(n925), .CK(i_clk), .RN(n470), .Q(n1649), .QN(n860)
         );
  DFFRX1 \LO_r_reg[4]  ( .D(n926), .CK(i_clk), .RN(n470), .Q(n1648), .QN(n859)
         );
  DFFRX1 \LO_r_reg[3]  ( .D(n927), .CK(i_clk), .RN(n470), .Q(n1647), .QN(n858)
         );
  DFFRX1 \LO_r_reg[2]  ( .D(n930), .CK(i_clk), .RN(n470), .Q(n1646), .QN(n855)
         );
  DFFRX1 \LO_r_reg[9]  ( .D(n921), .CK(i_clk), .RN(n470), .Q(n1653), .QN(n864)
         );
  DFFRX1 \HI_r_reg[9]  ( .D(n965), .CK(i_clk), .RN(n471), .Q(n1673), .QN(n831)
         );
  DFFRX1 \LO_r_reg[10]  ( .D(n961), .CK(i_clk), .RN(n470), .Q(n1654), .QN(n834) );
  DFFRX1 \HI_r_reg[10]  ( .D(n1286), .CK(i_clk), .RN(n471), .Q(n1674), .QN(
        n801) );
  DFFRX1 \LO_r_reg[11]  ( .D(n959), .CK(i_clk), .RN(n470), .Q(n1655), .QN(n835) );
  DFFRX1 \HI_r_reg[11]  ( .D(n1285), .CK(i_clk), .RN(n471), .Q(n1675), .QN(
        n802) );
  DFFRX1 \LO_r_reg[12]  ( .D(n957), .CK(i_clk), .RN(n470), .Q(n1656), .QN(n836) );
  DFFRX1 \HI_r_reg[12]  ( .D(n1284), .CK(i_clk), .RN(n471), .Q(n1676), .QN(
        n803) );
  DFFRX1 \LO_r_reg[13]  ( .D(n955), .CK(i_clk), .RN(n470), .Q(n1657), .QN(n837) );
  DFFRX1 \HI_r_reg[13]  ( .D(n1283), .CK(i_clk), .RN(n471), .Q(n1677), .QN(
        n804) );
  DFFRX1 \LO_r_reg[14]  ( .D(n953), .CK(i_clk), .RN(n470), .Q(n1658), .QN(n838) );
  DFFRX1 \HI_r_reg[14]  ( .D(n1282), .CK(i_clk), .RN(n471), .Q(n1678), .QN(
        n805) );
  DFFRX1 \LO_r_reg[15]  ( .D(n946), .CK(i_clk), .RN(n470), .Q(n1659), .QN(n839) );
  DFFRX1 \HI_r_reg[15]  ( .D(n1015), .CK(i_clk), .RN(n471), .Q(n1679), .QN(
        n806) );
  DFFRX1 \LO_r_reg[16]  ( .D(n945), .CK(i_clk), .RN(n470), .Q(n1660), .QN(n840) );
  DFFRX1 \HI_r_reg[16]  ( .D(n1013), .CK(i_clk), .RN(n471), .Q(n1680), .QN(
        n807) );
  DFFRX1 \LO_r_reg[17]  ( .D(n944), .CK(i_clk), .RN(n470), .Q(n1661), .QN(n841) );
  DFFRX1 \HI_r_reg[17]  ( .D(n1011), .CK(i_clk), .RN(n471), .Q(n1681), .QN(
        n808) );
  DFFRX1 \LO_r_reg[18]  ( .D(n943), .CK(i_clk), .RN(n470), .Q(n1662), .QN(n842) );
  DFFRX1 \HI_r_reg[18]  ( .D(n1009), .CK(i_clk), .RN(n471), .Q(n1682), .QN(
        n809) );
  DFFRX1 \LO_r_reg[19]  ( .D(n942), .CK(i_clk), .RN(n470), .Q(n1663), .QN(n843) );
  DFFRX1 \HI_r_reg[19]  ( .D(n1007), .CK(i_clk), .RN(n471), .Q(n1683), .QN(
        n810) );
  DFFRX2 \RegRd_memwb_r_reg[0]  ( .D(n1238), .CK(i_clk), .RN(n466), .Q(
        RegRd_memwb_r[0]), .QN(n1088) );
  DFFRX2 \RegRd_memwb_r_reg[4]  ( .D(n1236), .CK(i_clk), .RN(n460), .Q(
        RegRd_memwb_r[4]), .QN(n1086) );
  DFFRX2 \inst_r_reg[30]  ( .D(inst_w[30]), .CK(i_clk), .RN(n467), .Q(
        inst_r[30]), .QN(n913) );
  DFFRX2 \PC_r_reg[2]  ( .D(PC_w[2]), .CK(i_clk), .RN(n469), .Q(ICACHE_addr[0]) );
  DFFRX2 \PC_r_reg[4]  ( .D(PC_w[4]), .CK(i_clk), .RN(n469), .Q(ICACHE_addr[2]) );
  DFFRX2 \PC_r_reg[5]  ( .D(PC_w[5]), .CK(i_clk), .RN(n469), .Q(ICACHE_addr[3]) );
  OAI22X2 U40 ( .A0(n204), .A1(n1551), .B0(n1528), .B1(n207), .Y(ALUin2[2]) );
  OAI22X2 U41 ( .A0(n204), .A1(n1553), .B0(n456), .B1(n207), .Y(ALUin2[31]) );
  OAI22X2 U42 ( .A0(n204), .A1(n1554), .B0(n1472), .B1(n205), .Y(ALUin2[30])
         );
  OAI22X2 U43 ( .A0(n204), .A1(n1558), .B0(n1480), .B1(n44), .Y(ALUin2[26]) );
  OAI22X2 U44 ( .A0(n204), .A1(n1560), .B0(n1484), .B1(n44), .Y(ALUin2[24]) );
  OAI22X2 U45 ( .A0(n204), .A1(n1562), .B0(n1488), .B1(n206), .Y(ALUin2[22])
         );
  OAI22X2 U46 ( .A0(n204), .A1(n1564), .B0(n1492), .B1(n207), .Y(ALUin2[20])
         );
  OAI22X2 U47 ( .A0(n203), .A1(n1566), .B0(n1496), .B1(n206), .Y(ALUin2[18])
         );
  OAI22X2 U48 ( .A0(n203), .A1(n1567), .B0(n1498), .B1(n206), .Y(ALUin2[17])
         );
  OAI22X2 U49 ( .A0(n203), .A1(n1568), .B0(n1500), .B1(n205), .Y(ALUin2[16])
         );
  OAI22X2 U50 ( .A0(n203), .A1(n1571), .B0(n1504), .B1(n205), .Y(ALUin2[14])
         );
  OAI22X2 U51 ( .A0(n203), .A1(n1546), .B0(n1520), .B1(n206), .Y(ALUin2[6]) );
  CLKBUFX6 U52 ( .A(n476), .Y(n474) );
  CLKBUFX6 U53 ( .A(n476), .Y(n473) );
  CLKBUFX6 U54 ( .A(n478), .Y(n467) );
  CLKBUFX6 U55 ( .A(n479), .Y(n466) );
  CLKBUFX6 U56 ( .A(n477), .Y(n472) );
  CLKBUFX6 U57 ( .A(n479), .Y(n464) );
  CLKBUFX6 U58 ( .A(n480), .Y(n462) );
  CLKBUFX6 U59 ( .A(n480), .Y(n460) );
  CLKBUFX6 U60 ( .A(n478), .Y(n469) );
  AND2X2 U61 ( .A(n237), .B(n571), .Y(n42) );
  CLKBUFX2 U62 ( .A(n260), .Y(n263) );
  INVXL U63 ( .A(n1083), .Y(n70) );
  INVXL U64 ( .A(n1080), .Y(n71) );
  INVX3 U65 ( .A(n914), .Y(n72) );
  CLKINVX1 U66 ( .A(n1077), .Y(n73) );
  INVX16 U67 ( .A(n1096), .Y(DCACHE_wen) );
  CLKINVX1 U68 ( .A(n140), .Y(n75) );
  INVX16 U69 ( .A(n75), .Y(DCACHE_addr[1]) );
  CLKINVX1 U70 ( .A(n183), .Y(n77) );
  INVX16 U71 ( .A(n77), .Y(DCACHE_addr[0]) );
  CLKINVX1 U72 ( .A(n141), .Y(n79) );
  INVX16 U73 ( .A(n79), .Y(DCACHE_addr[3]) );
  CLKINVX1 U74 ( .A(n184), .Y(n81) );
  INVX16 U75 ( .A(n81), .Y(DCACHE_addr[2]) );
  CLKINVX1 U76 ( .A(n133), .Y(n83) );
  INVX16 U77 ( .A(n83), .Y(DCACHE_addr[29]) );
  CLKINVX1 U78 ( .A(n192), .Y(n85) );
  INVX16 U79 ( .A(n85), .Y(DCACHE_addr[28]) );
  CLKINVX1 U80 ( .A(n146), .Y(n87) );
  INVX16 U81 ( .A(n87), .Y(DCACHE_addr[27]) );
  CLKINVX1 U82 ( .A(n194), .Y(n89) );
  INVX16 U83 ( .A(n89), .Y(DCACHE_addr[26]) );
  CLKINVX1 U84 ( .A(n148), .Y(n91) );
  INVX16 U85 ( .A(n91), .Y(DCACHE_addr[25]) );
  CLKINVX1 U86 ( .A(n138), .Y(n93) );
  INVX16 U87 ( .A(n93), .Y(DCACHE_addr[24]) );
  CLKINVX1 U88 ( .A(n145), .Y(n95) );
  INVX16 U89 ( .A(n95), .Y(DCACHE_addr[23]) );
  CLKINVX1 U90 ( .A(n187), .Y(n97) );
  INVX16 U91 ( .A(n97), .Y(DCACHE_addr[22]) );
  CLKINVX1 U92 ( .A(n190), .Y(n99) );
  INVX16 U93 ( .A(n99), .Y(DCACHE_addr[21]) );
  CLKINVX1 U94 ( .A(n186), .Y(n101) );
  INVX16 U95 ( .A(n101), .Y(DCACHE_addr[20]) );
  CLKINVX1 U96 ( .A(n142), .Y(n103) );
  INVX16 U97 ( .A(n103), .Y(DCACHE_addr[19]) );
  CLKINVX1 U98 ( .A(n134), .Y(n105) );
  INVX16 U99 ( .A(n105), .Y(DCACHE_addr[18]) );
  CLKINVX1 U100 ( .A(n136), .Y(n107) );
  INVX16 U101 ( .A(n107), .Y(DCACHE_addr[17]) );
  CLKINVX1 U102 ( .A(n195), .Y(n109) );
  INVX16 U103 ( .A(n109), .Y(DCACHE_addr[16]) );
  CLKINVX1 U104 ( .A(n149), .Y(n111) );
  INVX16 U105 ( .A(n111), .Y(DCACHE_addr[15]) );
  CLKINVX1 U106 ( .A(n193), .Y(n113) );
  INVX16 U107 ( .A(n113), .Y(DCACHE_addr[14]) );
  CLKINVX1 U108 ( .A(n147), .Y(n115) );
  INVX16 U109 ( .A(n115), .Y(DCACHE_addr[13]) );
  CLKINVX1 U110 ( .A(n137), .Y(n117) );
  INVX16 U111 ( .A(n117), .Y(DCACHE_addr[12]) );
  CLKINVX1 U112 ( .A(n188), .Y(n119) );
  INVX16 U113 ( .A(n119), .Y(DCACHE_addr[11]) );
  CLKINVX1 U114 ( .A(n139), .Y(n121) );
  INVX16 U115 ( .A(n121), .Y(DCACHE_addr[10]) );
  CLKINVX1 U116 ( .A(n143), .Y(n123) );
  INVX16 U117 ( .A(n123), .Y(DCACHE_addr[9]) );
  CLKINVX1 U118 ( .A(n185), .Y(n125) );
  INVX16 U119 ( .A(n125), .Y(DCACHE_addr[8]) );
  CLKINVX1 U120 ( .A(n135), .Y(n127) );
  INVX16 U121 ( .A(n127), .Y(DCACHE_addr[7]) );
  CLKINVX1 U122 ( .A(n191), .Y(n129) );
  INVX16 U123 ( .A(n129), .Y(DCACHE_addr[6]) );
  CLKINVX1 U124 ( .A(n144), .Y(n131) );
  INVX16 U125 ( .A(n131), .Y(DCACHE_addr[5]) );
  BUFX12 U126 ( .A(n1684), .Y(DCACHE_addr[4]) );
  BUFX12 U127 ( .A(n1715), .Y(DCACHE_wdata[1]) );
  BUFX12 U128 ( .A(n1714), .Y(DCACHE_wdata[2]) );
  BUFX12 U129 ( .A(n1713), .Y(DCACHE_wdata[3]) );
  BUFX12 U130 ( .A(n1712), .Y(DCACHE_wdata[4]) );
  BUFX12 U131 ( .A(n1711), .Y(DCACHE_wdata[5]) );
  BUFX12 U132 ( .A(n1710), .Y(DCACHE_wdata[6]) );
  BUFX12 U133 ( .A(n1709), .Y(DCACHE_wdata[7]) );
  BUFX12 U134 ( .A(n1708), .Y(DCACHE_wdata[8]) );
  BUFX12 U135 ( .A(n1707), .Y(DCACHE_wdata[9]) );
  BUFX12 U136 ( .A(n1706), .Y(DCACHE_wdata[10]) );
  BUFX12 U137 ( .A(n1705), .Y(DCACHE_wdata[11]) );
  BUFX12 U138 ( .A(n1704), .Y(DCACHE_wdata[12]) );
  BUFX12 U139 ( .A(n1703), .Y(DCACHE_wdata[13]) );
  BUFX12 U140 ( .A(n1702), .Y(DCACHE_wdata[14]) );
  BUFX12 U141 ( .A(n1701), .Y(DCACHE_wdata[15]) );
  BUFX12 U142 ( .A(n1700), .Y(DCACHE_wdata[16]) );
  BUFX12 U143 ( .A(n1699), .Y(DCACHE_wdata[17]) );
  BUFX12 U144 ( .A(n1698), .Y(DCACHE_wdata[18]) );
  BUFX12 U145 ( .A(n1697), .Y(DCACHE_wdata[19]) );
  BUFX12 U146 ( .A(n1696), .Y(DCACHE_wdata[20]) );
  BUFX12 U147 ( .A(n1695), .Y(DCACHE_wdata[21]) );
  BUFX12 U148 ( .A(n1694), .Y(DCACHE_wdata[22]) );
  BUFX12 U149 ( .A(n1693), .Y(DCACHE_wdata[23]) );
  BUFX12 U150 ( .A(n1692), .Y(DCACHE_wdata[24]) );
  BUFX12 U151 ( .A(n1691), .Y(DCACHE_wdata[25]) );
  BUFX12 U152 ( .A(n1690), .Y(DCACHE_wdata[26]) );
  BUFX12 U153 ( .A(n1689), .Y(DCACHE_wdata[27]) );
  BUFX12 U154 ( .A(n1688), .Y(DCACHE_wdata[28]) );
  BUFX12 U155 ( .A(n1687), .Y(DCACHE_wdata[29]) );
  BUFX12 U156 ( .A(n1685), .Y(DCACHE_wdata[31]) );
  BUFX12 U157 ( .A(n1686), .Y(DCACHE_wdata[30]) );
  BUFX12 U158 ( .A(n1716), .Y(DCACHE_wdata[0]) );
  BUFX4 U159 ( .A(n480), .Y(n458) );
  NAND2X1 U160 ( .A(n570), .B(n238), .Y(n507) );
  NAND2X1 U161 ( .A(n219), .B(n222), .Y(n725) );
  NAND2X1 U162 ( .A(n227), .B(n229), .Y(n722) );
  CLKINVX1 U163 ( .A(n508), .Y(n237) );
  NAND2BX1 U164 ( .AN(forwardB[1]), .B(n199), .Y(n790) );
  NAND2X1 U165 ( .A(forwardB[1]), .B(n199), .Y(n792) );
  NAND2BX1 U166 ( .AN(forwardA[1]), .B(n201), .Y(n395) );
  NAND2X1 U167 ( .A(forwardA[1]), .B(n201), .Y(n394) );
  AND4X1 U168 ( .A(JumpR), .B(PCSrc), .C(n238), .D(n693), .Y(n501) );
  AND4X1 U169 ( .A(n686), .B(ICACHE_rdata[28]), .C(n238), .D(n700), .Y(n509)
         );
  NAND2BX1 U170 ( .AN(ForwardJB[1]), .B(ForwardJB[0]), .Y(n720) );
  NAND2BX1 U171 ( .AN(ForwardJA[1]), .B(ForwardJA[0]), .Y(n723) );
  NAND2BX1 U172 ( .AN(ForwardJB[0]), .B(ForwardJB[1]), .Y(n721) );
  NAND2BX1 U173 ( .AN(ForwardJA[0]), .B(ForwardJA[1]), .Y(n724) );
  CLKINVX1 U174 ( .A(readreg2_forward[31]), .Y(n456) );
  CLKINVX1 U175 ( .A(forwardB[0]), .Y(n1534) );
  OAI222X1 U176 ( .A0(n1580), .A1(n216), .B0(n199), .B1(n396), .C0(n1429), 
        .C1(n214), .Y(readreg2_forward[0]) );
  OAI222X1 U177 ( .A0(n1581), .A1(n216), .B0(n199), .B1(n420), .C0(n1428), 
        .C1(n214), .Y(readreg2_forward[1]) );
  CLKBUFX3 U178 ( .A(n1105), .Y(n212) );
  OAI2BB2X1 U179 ( .B0(n211), .B1(n1137), .A0N(n212), .A1N(n1102), .Y(n447) );
  CLKINVX1 U180 ( .A(forwardA[0]), .Y(n1535) );
  OAI222X1 U181 ( .A0(n1427), .A1(n249), .B0(n1614), .B1(n247), .C0(n443), 
        .C1(n201), .Y(readreg1_forward[2]) );
  OAI222X1 U182 ( .A0(n1428), .A1(n248), .B0(n1613), .B1(n246), .C0(n420), 
        .C1(n202), .Y(readreg1_forward[1]) );
  OAI222X1 U183 ( .A0(n1429), .A1(n248), .B0(n1612), .B1(n246), .C0(n396), 
        .C1(n201), .Y(readreg1_forward[0]) );
  OAI222X1 U184 ( .A0(n1582), .A1(n215), .B0(n200), .B1(n443), .C0(n1427), 
        .C1(n213), .Y(readreg2_forward[2]) );
  OAI222X1 U185 ( .A0(n1583), .A1(n215), .B0(n200), .B1(n450), .C0(n1426), 
        .C1(n213), .Y(readreg2_forward[3]) );
  OAI222X1 U186 ( .A0(n1584), .A1(n215), .B0(n200), .B1(n453), .C0(n1425), 
        .C1(n213), .Y(readreg2_forward[4]) );
  OAI222X1 U187 ( .A0(n1585), .A1(n215), .B0(n200), .B1(n455), .C0(n1424), 
        .C1(n213), .Y(readreg2_forward[5]) );
  OAI2BB2X1 U188 ( .B0(n211), .B1(n1109), .A0N(n212), .A1N(n1071), .Y(n450) );
  OAI2BB2X1 U189 ( .B0(n210), .B1(n1106), .A0N(n209), .A1N(n1100), .Y(n396) );
  OAI2BB2X1 U190 ( .B0(n210), .B1(n1108), .A0N(n212), .A1N(n1073), .Y(n443) );
  OAI2BB2X1 U191 ( .B0(n209), .B1(n1107), .A0N(n212), .A1N(n1075), .Y(n420) );
  OAI222X1 U192 ( .A0(n1425), .A1(n249), .B0(n1616), .B1(n247), .C0(n453), 
        .C1(n201), .Y(readreg1_forward[4]) );
  OAI222X1 U193 ( .A0(n1426), .A1(n249), .B0(n1615), .B1(n247), .C0(n450), 
        .C1(n202), .Y(readreg1_forward[3]) );
  OAI222X1 U194 ( .A0(n1588), .A1(n215), .B0(n199), .B1(n461), .C0(n1421), 
        .C1(n213), .Y(readreg2_forward[8]) );
  OAI222X1 U195 ( .A0(n1586), .A1(n215), .B0(n200), .B1(n457), .C0(n1423), 
        .C1(n213), .Y(readreg2_forward[6]) );
  OAI222X1 U196 ( .A0(n1587), .A1(n215), .B0(n199), .B1(n459), .C0(n1422), 
        .C1(n213), .Y(readreg2_forward[7]) );
  OAI2BB2X1 U197 ( .B0(n211), .B1(n1112), .A0N(n212), .A1N(n1065), .Y(n457) );
  OAI2BB2X1 U198 ( .B0(n211), .B1(n1111), .A0N(n212), .A1N(n1067), .Y(n455) );
  OAI2BB2X1 U199 ( .B0(n211), .B1(n1110), .A0N(n212), .A1N(n1069), .Y(n453) );
  NAND3BX1 U200 ( .AN(n832), .B(n903), .C(n799), .Y(n393) );
  NAND3X1 U201 ( .A(n832), .B(n903), .C(n799), .Y(n390) );
  OR2X1 U202 ( .A(n799), .B(n43), .Y(n388) );
  OAI222X1 U203 ( .A0(n1421), .A1(n249), .B0(n1620), .B1(n247), .C0(n461), 
        .C1(n201), .Y(readreg1_forward[8]) );
  OAI222X1 U204 ( .A0(n1423), .A1(n249), .B0(n1618), .B1(n247), .C0(n457), 
        .C1(n201), .Y(readreg1_forward[6]) );
  OAI222X1 U205 ( .A0(n1422), .A1(n249), .B0(n1619), .B1(n247), .C0(n459), 
        .C1(n201), .Y(readreg1_forward[7]) );
  OAI222X1 U206 ( .A0(n1424), .A1(n249), .B0(n1617), .B1(n247), .C0(n455), 
        .C1(n201), .Y(readreg1_forward[5]) );
  OAI222X1 U207 ( .A0(n1589), .A1(n215), .B0(n463), .B1(n199), .C0(n1420), 
        .C1(n213), .Y(readreg2_forward[9]) );
  OAI222X1 U208 ( .A0(n1590), .A1(n216), .B0(n199), .B1(n399), .C0(n1419), 
        .C1(n214), .Y(readreg2_forward[10]) );
  OAI222X1 U209 ( .A0(n1591), .A1(n216), .B0(n199), .B1(n401), .C0(n1418), 
        .C1(n214), .Y(readreg2_forward[11]) );
  OAI2BB2X1 U210 ( .B0(n211), .B1(n1114), .A0N(n209), .A1N(n1061), .Y(n461) );
  OAI2BB2X1 U211 ( .B0(n211), .B1(n1113), .A0N(n212), .A1N(n1063), .Y(n459) );
  OAI2BB2X1 U212 ( .B0(n211), .B1(n1115), .A0N(n210), .A1N(n1059), .Y(n463) );
  OAI222X1 U213 ( .A0(n1420), .A1(n249), .B0(n1621), .B1(n247), .C0(n463), 
        .C1(n201), .Y(readreg1_forward[9]) );
  OAI222X1 U214 ( .A0(n1419), .A1(n248), .B0(n1622), .B1(n246), .C0(n399), 
        .C1(n202), .Y(readreg1_forward[10]) );
  OAI222X1 U215 ( .A0(n1418), .A1(n248), .B0(n1623), .B1(n246), .C0(n401), 
        .C1(n202), .Y(readreg1_forward[11]) );
  OAI222X1 U216 ( .A0(n1592), .A1(n216), .B0(n199), .B1(n403), .C0(n1417), 
        .C1(n214), .Y(readreg2_forward[12]) );
  OAI222X1 U217 ( .A0(n1593), .A1(n216), .B0(n199), .B1(n405), .C0(n1416), 
        .C1(n214), .Y(readreg2_forward[13]) );
  OAI222X1 U218 ( .A0(n1594), .A1(n216), .B0(n199), .B1(n407), .C0(n1415), 
        .C1(n214), .Y(readreg2_forward[14]) );
  OAI2BB2X1 U219 ( .B0(n209), .B1(n1119), .A0N(n212), .A1N(n1051), .Y(n405) );
  OAI2BB2X1 U220 ( .B0(n209), .B1(n1116), .A0N(n209), .A1N(n1057), .Y(n399) );
  OAI2BB2X1 U221 ( .B0(n209), .B1(n1117), .A0N(n210), .A1N(n1055), .Y(n401) );
  OAI2BB2X1 U222 ( .B0(n209), .B1(n1118), .A0N(n212), .A1N(n1053), .Y(n403) );
  OAI222X1 U223 ( .A0(n1416), .A1(n248), .B0(n1625), .B1(n246), .C0(n405), 
        .C1(n202), .Y(readreg1_forward[13]) );
  OAI222X1 U224 ( .A0(n1415), .A1(n248), .B0(n1626), .B1(n246), .C0(n407), 
        .C1(n201), .Y(readreg1_forward[14]) );
  OAI222X1 U225 ( .A0(n1414), .A1(n248), .B0(n1627), .B1(n246), .C0(n409), 
        .C1(n202), .Y(readreg1_forward[15]) );
  OAI222X1 U226 ( .A0(n1417), .A1(n248), .B0(n1624), .B1(n246), .C0(n403), 
        .C1(n202), .Y(readreg1_forward[12]) );
  OAI222X1 U227 ( .A0(n1596), .A1(n215), .B0(n199), .B1(n411), .C0(n1413), 
        .C1(n214), .Y(readreg2_forward[16]) );
  OAI222X1 U228 ( .A0(n1597), .A1(n216), .B0(n199), .B1(n413), .C0(n1412), 
        .C1(n214), .Y(readreg2_forward[17]) );
  OAI222X1 U229 ( .A0(n1595), .A1(n216), .B0(n200), .B1(n409), .C0(n1414), 
        .C1(n214), .Y(readreg2_forward[15]) );
  OAI2BB2X1 U230 ( .B0(n209), .B1(n1120), .A0N(n212), .A1N(n1049), .Y(n407) );
  OAI2BB2X1 U231 ( .B0(n209), .B1(n1121), .A0N(n212), .A1N(n1047), .Y(n409) );
  OAI2BB2X1 U232 ( .B0(n209), .B1(n1122), .A0N(n212), .A1N(n1045), .Y(n411) );
  OAI222X1 U233 ( .A0(n1412), .A1(n248), .B0(n1629), .B1(n246), .C0(n413), 
        .C1(n202), .Y(readreg1_forward[17]) );
  OAI222X1 U234 ( .A0(n1411), .A1(n248), .B0(n1630), .B1(n246), .C0(n415), 
        .C1(n202), .Y(readreg1_forward[18]) );
  OAI222X1 U235 ( .A0(n1413), .A1(n248), .B0(n1628), .B1(n246), .C0(n411), 
        .C1(n202), .Y(readreg1_forward[16]) );
  OAI222X1 U236 ( .A0(n1598), .A1(n216), .B0(n199), .B1(n415), .C0(n1411), 
        .C1(n214), .Y(readreg2_forward[18]) );
  OAI222X1 U237 ( .A0(n1599), .A1(n216), .B0(n199), .B1(n417), .C0(n1410), 
        .C1(n214), .Y(readreg2_forward[19]) );
  OAI222X1 U238 ( .A0(n1600), .A1(n216), .B0(n200), .B1(n422), .C0(n1409), 
        .C1(n214), .Y(readreg2_forward[20]) );
  OAI222X1 U239 ( .A0(n1601), .A1(n216), .B0(n200), .B1(n424), .C0(n1408), 
        .C1(n214), .Y(readreg2_forward[21]) );
  OAI2BB2X1 U240 ( .B0(n209), .B1(n1123), .A0N(n212), .A1N(n1043), .Y(n413) );
  OAI2BB2X1 U241 ( .B0(n209), .B1(n1124), .A0N(n209), .A1N(n1041), .Y(n415) );
  OAI2BB2X1 U242 ( .B0(n209), .B1(n1125), .A0N(n212), .A1N(n1039), .Y(n417) );
  OAI222X1 U243 ( .A0(n1410), .A1(n248), .B0(n1631), .B1(n246), .C0(n417), 
        .C1(n202), .Y(readreg1_forward[19]) );
  OAI222X1 U244 ( .A0(n1409), .A1(n249), .B0(n1632), .B1(n247), .C0(n422), 
        .C1(n202), .Y(readreg1_forward[20]) );
  OAI222X1 U245 ( .A0(n1408), .A1(n249), .B0(n1633), .B1(n247), .C0(n424), 
        .C1(n202), .Y(readreg1_forward[21]) );
  OAI222X1 U246 ( .A0(n1602), .A1(n216), .B0(n200), .B1(n426), .C0(n1407), 
        .C1(n214), .Y(readreg2_forward[22]) );
  OAI222X1 U247 ( .A0(n1603), .A1(n216), .B0(n200), .B1(n428), .C0(n1406), 
        .C1(n214), .Y(readreg2_forward[23]) );
  OAI222X1 U248 ( .A0(n1604), .A1(n216), .B0(n200), .B1(n430), .C0(n1405), 
        .C1(n214), .Y(readreg2_forward[24]) );
  OAI222XL U249 ( .A0(n1428), .A1(n222), .B0(n420), .B1(n219), .C0(n1466), 
        .C1(n218), .Y(n625) );
  OAI222XL U250 ( .A0(n1410), .A1(n222), .B0(n417), .B1(n219), .C0(n1314), 
        .C1(n217), .Y(n629) );
  OAI222XL U251 ( .A0(n1414), .A1(n222), .B0(n409), .B1(n219), .C0(n1322), 
        .C1(n217), .Y(n653) );
  OAI222XL U252 ( .A0(n1415), .A1(n222), .B0(n407), .B1(n219), .C0(n1324), 
        .C1(n217), .Y(n659) );
  OAI222XL U253 ( .A0(n1416), .A1(n222), .B0(n405), .B1(n219), .C0(n1326), 
        .C1(n217), .Y(n665) );
  OAI222XL U254 ( .A0(n1417), .A1(n222), .B0(n403), .B1(n219), .C0(n1328), 
        .C1(n218), .Y(n671) );
  OAI222XL U255 ( .A0(n1419), .A1(n222), .B0(n399), .B1(n219), .C0(n1332), 
        .C1(n217), .Y(n683) );
  OAI222XL U256 ( .A0(n1420), .A1(n222), .B0(n463), .B1(n219), .C0(n1334), 
        .C1(n217), .Y(n502) );
  OAI222XL U257 ( .A0(n1421), .A1(n222), .B0(n461), .B1(n219), .C0(n1336), 
        .C1(n217), .Y(n514) );
  OAI222XL U258 ( .A0(n1422), .A1(n222), .B0(n459), .B1(n219), .C0(n1338), 
        .C1(n217), .Y(n520) );
  OAI222XL U259 ( .A0(n1423), .A1(n222), .B0(n457), .B1(n219), .C0(n1340), 
        .C1(n217), .Y(n526) );
  OAI222XL U260 ( .A0(n1424), .A1(n222), .B0(n455), .B1(n219), .C0(n1342), 
        .C1(n217), .Y(n532) );
  OAI222XL U261 ( .A0(n1425), .A1(n222), .B0(n453), .B1(n219), .C0(n1344), 
        .C1(n217), .Y(n538) );
  OAI222XL U262 ( .A0(n1398), .A1(n224), .B0(n447), .B1(n220), .C0(n1290), 
        .C1(n218), .Y(n551) );
  OAI222XL U263 ( .A0(n1399), .A1(n224), .B0(n445), .B1(n220), .C0(n1292), 
        .C1(n218), .Y(n555) );
  OAI222XL U264 ( .A0(n1400), .A1(n224), .B0(n440), .B1(n220), .C0(n1294), 
        .C1(n218), .Y(n565) );
  OAI222XL U265 ( .A0(n1401), .A1(n224), .B0(n438), .B1(n220), .C0(n1296), 
        .C1(n218), .Y(n569) );
  OAI222XL U266 ( .A0(n1402), .A1(n224), .B0(n436), .B1(n220), .C0(n1298), 
        .C1(n218), .Y(n576) );
  OAI222XL U267 ( .A0(n1403), .A1(n224), .B0(n434), .B1(n220), .C0(n1300), 
        .C1(n218), .Y(n582) );
  OAI222XL U268 ( .A0(n1404), .A1(n224), .B0(n432), .B1(n220), .C0(n1302), 
        .C1(n218), .Y(n588) );
  OAI222XL U269 ( .A0(n1405), .A1(n224), .B0(n430), .B1(n220), .C0(n1304), 
        .C1(n218), .Y(n594) );
  OAI222XL U270 ( .A0(n1406), .A1(n224), .B0(n428), .B1(n220), .C0(n1306), 
        .C1(n218), .Y(n600) );
  OAI222XL U271 ( .A0(n1407), .A1(n224), .B0(n426), .B1(n220), .C0(n1308), 
        .C1(n217), .Y(n606) );
  OAI222XL U272 ( .A0(n1408), .A1(n224), .B0(n424), .B1(n220), .C0(n1310), 
        .C1(n725), .Y(n612) );
  OAI222XL U273 ( .A0(n1409), .A1(n224), .B0(n422), .B1(n220), .C0(n1312), 
        .C1(n218), .Y(n618) );
  OAI222XL U274 ( .A0(n1418), .A1(n224), .B0(n401), .B1(n220), .C0(n1330), 
        .C1(n217), .Y(n677) );
  OAI222XL U275 ( .A0(n1426), .A1(n224), .B0(n450), .B1(n220), .C0(n1462), 
        .C1(n218), .Y(n544) );
  OAI222XL U276 ( .A0(n1427), .A1(n222), .B0(n443), .B1(n220), .C0(n1464), 
        .C1(n218), .Y(n559) );
  OAI222XL U277 ( .A0(n1468), .A1(n217), .B0(n1429), .B1(n224), .C0(n396), 
        .C1(n219), .Y(n692) );
  OAI222XL U278 ( .A0(n1411), .A1(n224), .B0(n415), .B1(n220), .C0(n1316), 
        .C1(n725), .Y(n635) );
  OAI222XL U279 ( .A0(n1412), .A1(n224), .B0(n413), .B1(n220), .C0(n1318), 
        .C1(n725), .Y(n641) );
  OAI222XL U280 ( .A0(n1413), .A1(n224), .B0(n411), .B1(n220), .C0(n1320), 
        .C1(n725), .Y(n647) );
  OAI2BB2X1 U281 ( .B0(n209), .B1(n1126), .A0N(n212), .A1N(n1037), .Y(n422) );
  OAI2BB2X1 U282 ( .B0(n210), .B1(n1127), .A0N(n212), .A1N(n1035), .Y(n424) );
  OAI2BB2X1 U283 ( .B0(n210), .B1(n1128), .A0N(n212), .A1N(n1033), .Y(n426) );
  OAI21XL U284 ( .A0(n693), .A1(n1289), .B0(n695), .Y(n571) );
  NAND2X1 U285 ( .A(n1396), .B(n307), .Y(n223) );
  OR2X1 U286 ( .A(n1396), .B(n345), .Y(n221) );
  OAI222X1 U287 ( .A0(n1405), .A1(n249), .B0(n1636), .B1(n247), .C0(n430), 
        .C1(n202), .Y(readreg1_forward[24]) );
  OAI222X1 U288 ( .A0(n1407), .A1(n249), .B0(n1634), .B1(n247), .C0(n426), 
        .C1(n202), .Y(readreg1_forward[22]) );
  OAI222X1 U289 ( .A0(n1406), .A1(n249), .B0(n1635), .B1(n247), .C0(n428), 
        .C1(n202), .Y(readreg1_forward[23]) );
  OAI222X1 U290 ( .A0(n1404), .A1(n249), .B0(n1637), .B1(n247), .C0(n432), 
        .C1(n202), .Y(readreg1_forward[25]) );
  OAI222X1 U291 ( .A0(n1605), .A1(n216), .B0(n200), .B1(n432), .C0(n1404), 
        .C1(n214), .Y(readreg2_forward[25]) );
  OAI222X1 U292 ( .A0(n1606), .A1(n216), .B0(n200), .B1(n434), .C0(n1403), 
        .C1(n214), .Y(readreg2_forward[26]) );
  OAI222X1 U293 ( .A0(n1607), .A1(n216), .B0(n200), .B1(n436), .C0(n1402), 
        .C1(n213), .Y(readreg2_forward[27]) );
  OAI2BB2X1 U294 ( .B0(n210), .B1(n1129), .A0N(n211), .A1N(n1031), .Y(n428) );
  OAI2BB2X1 U295 ( .B0(n210), .B1(n1130), .A0N(n212), .A1N(n1029), .Y(n430) );
  OAI2BB2X1 U296 ( .B0(n210), .B1(n1131), .A0N(n211), .A1N(n1027), .Y(n432) );
  OAI2BB2X1 U297 ( .B0(n210), .B1(n1132), .A0N(n211), .A1N(n1025), .Y(n434) );
  OAI2BB2X1 U298 ( .B0(n210), .B1(n1133), .A0N(n212), .A1N(n1023), .Y(n436) );
  OAI2BB2X1 U299 ( .B0(n210), .B1(n1134), .A0N(n211), .A1N(n1021), .Y(n438) );
  OAI2BB2X1 U300 ( .B0(n210), .B1(n1135), .A0N(n211), .A1N(n1019), .Y(n440) );
  OAI2BB2X1 U301 ( .B0(n210), .B1(n1136), .A0N(n211), .A1N(n1017), .Y(n445) );
  CLKBUFX3 U302 ( .A(sign_ext_31), .Y(n198) );
  OAI222X1 U303 ( .A0(n1403), .A1(n249), .B0(n1638), .B1(n247), .C0(n434), 
        .C1(n202), .Y(readreg1_forward[26]) );
  OAI222X1 U304 ( .A0(n1402), .A1(n249), .B0(n1639), .B1(n247), .C0(n436), 
        .C1(n202), .Y(readreg1_forward[27]) );
  OAI222X1 U305 ( .A0(n1401), .A1(n249), .B0(n1640), .B1(n247), .C0(n438), 
        .C1(n201), .Y(readreg1_forward[28]) );
  OAI222X1 U306 ( .A0(n1400), .A1(n249), .B0(n1641), .B1(n247), .C0(n440), 
        .C1(n201), .Y(readreg1_forward[29]) );
  OAI222X1 U307 ( .A0(n1399), .A1(n248), .B0(n1642), .B1(n247), .C0(n445), 
        .C1(n201), .Y(readreg1_forward[30]) );
  OAI222X1 U308 ( .A0(n1398), .A1(n249), .B0(n1643), .B1(n246), .C0(n447), 
        .C1(n201), .Y(readreg1_forward[31]) );
  OAI222X1 U309 ( .A0(n1608), .A1(n215), .B0(n200), .B1(n438), .C0(n1401), 
        .C1(n213), .Y(readreg2_forward[28]) );
  OAI222X1 U310 ( .A0(n1609), .A1(n215), .B0(n200), .B1(n440), .C0(n1400), 
        .C1(n213), .Y(readreg2_forward[29]) );
  OAI222X1 U311 ( .A0(n1610), .A1(n215), .B0(n200), .B1(n445), .C0(n1399), 
        .C1(n213), .Y(readreg2_forward[30]) );
  AOI2BB1X1 U312 ( .A0N(n1397), .A1N(stall_div), .B0(n279), .Y(n260) );
  NOR2X1 U313 ( .A(n865), .B(stall_mul), .Y(n258) );
  INVX3 U314 ( .A(n389), .Y(n387) );
  INVX3 U315 ( .A(n397), .Y(n373) );
  INVX3 U316 ( .A(n406), .Y(n375) );
  INVX3 U317 ( .A(n402), .Y(n383) );
  INVX3 U318 ( .A(n404), .Y(n381) );
  INVX3 U319 ( .A(n400), .Y(n377) );
  INVX3 U320 ( .A(n408), .Y(n379) );
  INVX3 U321 ( .A(n389), .Y(n385) );
  CLKBUFX3 U322 ( .A(n429), .Y(n389) );
  CLKBUFX3 U323 ( .A(n429), .Y(n392) );
  CLKBUFX3 U324 ( .A(n392), .Y(n397) );
  CLKBUFX3 U325 ( .A(n414), .Y(n418) );
  CLKBUFX3 U326 ( .A(n410), .Y(n421) );
  CLKBUFX3 U327 ( .A(n427), .Y(n414) );
  CLKBUFX3 U328 ( .A(n414), .Y(n416) );
  CLKBUFX3 U329 ( .A(n427), .Y(n412) );
  CLKBUFX3 U330 ( .A(n433), .Y(n400) );
  CLKBUFX3 U331 ( .A(n433), .Y(n404) );
  CLKBUFX3 U332 ( .A(n433), .Y(n402) );
  CLKBUFX3 U333 ( .A(n433), .Y(n408) );
  CLKBUFX3 U334 ( .A(n433), .Y(n406) );
  CLKBUFX3 U335 ( .A(n392), .Y(n398) );
  CLKBUFX3 U336 ( .A(n427), .Y(n410) );
  CLKBUFX3 U337 ( .A(n507), .Y(n239) );
  CLKBUFX3 U338 ( .A(n510), .Y(n231) );
  CLKBUFX3 U339 ( .A(n510), .Y(n232) );
  CLKBUFX3 U340 ( .A(n431), .Y(n429) );
  INVX3 U341 ( .A(n355), .Y(n311) );
  INVX3 U342 ( .A(n317), .Y(n307) );
  INVX3 U343 ( .A(n367), .Y(n309) );
  INVX3 U344 ( .A(n355), .Y(n313) );
  CLKBUFX3 U345 ( .A(n410), .Y(n423) );
  CLKBUFX3 U346 ( .A(n722), .Y(n225) );
  CLKBUFX3 U347 ( .A(n725), .Y(n217) );
  CLKBUFX3 U348 ( .A(n725), .Y(n218) );
  INVX3 U349 ( .A(n357), .Y(n315) );
  CLKBUFX3 U350 ( .A(n722), .Y(n226) );
  CLKBUFX3 U351 ( .A(n435), .Y(n427) );
  CLKBUFX3 U352 ( .A(n398), .Y(n425) );
  INVX3 U353 ( .A(n355), .Y(n297) );
  INVX3 U354 ( .A(n359), .Y(n305) );
  INVX3 U355 ( .A(n359), .Y(n303) );
  INVX3 U356 ( .A(n357), .Y(n301) );
  INVX3 U357 ( .A(n355), .Y(n299) );
  CLKBUFX6 U358 ( .A(n477), .Y(n470) );
  CLKBUFX6 U359 ( .A(n477), .Y(n471) );
  CLKBUFX6 U360 ( .A(n479), .Y(n465) );
  CLKBUFX6 U361 ( .A(n478), .Y(n468) );
  CLKBUFX3 U362 ( .A(n476), .Y(n475) );
  CLKBUFX3 U363 ( .A(n444), .Y(n446) );
  CLKBUFX3 U364 ( .A(n13), .Y(n439) );
  CLKBUFX3 U365 ( .A(n13), .Y(n441) );
  CLKBUFX3 U366 ( .A(n13), .Y(n437) );
  INVX3 U367 ( .A(n237), .Y(n235) );
  CLKBUFX3 U368 ( .A(n361), .Y(n319) );
  INVX3 U369 ( .A(n42), .Y(n241) );
  INVX3 U370 ( .A(n42), .Y(n240) );
  CLKBUFX3 U371 ( .A(n503), .Y(n242) );
  CLKBUFX3 U372 ( .A(n503), .Y(n243) );
  CLKINVX1 U373 ( .A(n371), .Y(n431) );
  CLKBUFX3 U374 ( .A(n448), .Y(n451) );
  CLKBUFX3 U375 ( .A(n444), .Y(n448) );
  INVX3 U376 ( .A(n237), .Y(n236) );
  CLKBUFX3 U377 ( .A(n363), .Y(n317) );
  CLKBUFX3 U378 ( .A(n353), .Y(n345) );
  CLKBUFX3 U379 ( .A(n357), .Y(n337) );
  CLKBUFX3 U380 ( .A(n357), .Y(n335) );
  CLKBUFX3 U381 ( .A(n359), .Y(n333) );
  CLKBUFX3 U382 ( .A(n359), .Y(n331) );
  CLKBUFX3 U383 ( .A(n359), .Y(n329) );
  CLKBUFX3 U384 ( .A(n359), .Y(n327) );
  CLKBUFX3 U385 ( .A(n359), .Y(n325) );
  CLKBUFX3 U386 ( .A(n359), .Y(n323) );
  CLKBUFX3 U387 ( .A(n361), .Y(n321) );
  CLKINVX1 U388 ( .A(n371), .Y(n433) );
  CLKINVX1 U389 ( .A(n385), .Y(n435) );
  CLKBUFX3 U390 ( .A(n353), .Y(n347) );
  CLKBUFX3 U391 ( .A(n353), .Y(n349) );
  CLKBUFX3 U392 ( .A(n355), .Y(n343) );
  CLKBUFX3 U393 ( .A(n355), .Y(n341) );
  CLKBUFX3 U394 ( .A(n355), .Y(n339) );
  CLKBUFX3 U395 ( .A(n353), .Y(n351) );
  CLKBUFX3 U396 ( .A(rst_n), .Y(n480) );
  CLKBUFX3 U397 ( .A(rst_n), .Y(n477) );
  CLKBUFX3 U398 ( .A(n479), .Y(n476) );
  CLKBUFX3 U399 ( .A(n480), .Y(n478) );
  CLKBUFX3 U400 ( .A(rst_n), .Y(n479) );
  CLKBUFX3 U401 ( .A(n792), .Y(n213) );
  CLKBUFX3 U402 ( .A(n790), .Y(n216) );
  CLKBUFX3 U403 ( .A(n790), .Y(n215) );
  CLKBUFX3 U404 ( .A(n792), .Y(n214) );
  CLKBUFX3 U405 ( .A(n394), .Y(n248) );
  CLKBUFX3 U406 ( .A(n395), .Y(n246) );
  CLKBUFX3 U407 ( .A(n395), .Y(n247) );
  CLKBUFX3 U408 ( .A(n394), .Y(n249) );
  NOR3X1 U409 ( .A(n235), .B(PCSrc), .C(n1288), .Y(n510) );
  OAI22XL U410 ( .A0(n241), .A1(n602), .B0(n655), .B1(n239), .Y(n642) );
  OAI22XL U411 ( .A0(n241), .A1(n603), .B0(n656), .B1(n239), .Y(n648) );
  OAI22XL U412 ( .A0(n241), .A1(n608), .B0(n661), .B1(n239), .Y(n654) );
  OAI22XL U413 ( .A0(n241), .A1(n609), .B0(n662), .B1(n239), .Y(n660) );
  OAI22XL U414 ( .A0(n241), .A1(n614), .B0(n667), .B1(n239), .Y(n666) );
  OAI22XL U415 ( .A0(n241), .A1(n615), .B0(n668), .B1(n239), .Y(n672) );
  OAI22XL U416 ( .A0(n241), .A1(n620), .B0(n673), .B1(n507), .Y(n678) );
  OAI22XL U417 ( .A0(n241), .A1(n621), .B0(n674), .B1(n239), .Y(n684) );
  OAI22XL U418 ( .A0(n240), .A1(n624), .B0(n679), .B1(n507), .Y(n504) );
  OAI22XL U419 ( .A0(n240), .A1(n626), .B0(n680), .B1(n239), .Y(n515) );
  OAI22XL U420 ( .A0(n240), .A1(n631), .B0(n685), .B1(n507), .Y(n521) );
  OAI22XL U421 ( .A0(n240), .A1(n632), .B0(n688), .B1(n507), .Y(n527) );
  OAI22XL U422 ( .A0(n240), .A1(n637), .B0(n689), .B1(n239), .Y(n533) );
  OAI22XL U423 ( .A0(n240), .A1(n638), .B0(n694), .B1(n239), .Y(n539) );
  OAI22XL U424 ( .A0(n240), .A1(n643), .B0(n697), .B1(n239), .Y(n545) );
  OAI22XL U425 ( .A0(n240), .A1(n572), .B0(n789), .B1(n507), .Y(n577) );
  OAI22XL U426 ( .A0(n240), .A1(n573), .B0(n791), .B1(n507), .Y(n583) );
  OAI22XL U427 ( .A0(n240), .A1(n578), .B0(n915), .B1(n239), .Y(n589) );
  OAI22XL U428 ( .A0(n240), .A1(n579), .B0(n916), .B1(n239), .Y(n595) );
  OAI22XL U429 ( .A0(n241), .A1(n584), .B0(n917), .B1(n239), .Y(n601) );
  OAI22XL U430 ( .A0(n241), .A1(n585), .B0(n918), .B1(n239), .Y(n607) );
  OAI22XL U431 ( .A0(n241), .A1(n590), .B0(n919), .B1(n239), .Y(n613) );
  OAI22XL U432 ( .A0(n241), .A1(n591), .B0(n920), .B1(n239), .Y(n619) );
  OAI22XL U433 ( .A0(n241), .A1(n596), .B0(n649), .B1(n239), .Y(n630) );
  OAI22XL U434 ( .A0(n241), .A1(n597), .B0(n650), .B1(n239), .Y(n636) );
  INVX4 U435 ( .A(n208), .Y(n203) );
  INVX4 U436 ( .A(n206), .Y(n204) );
  CLKBUFX3 U437 ( .A(n208), .Y(n207) );
  CLKBUFX3 U438 ( .A(n208), .Y(n206) );
  CLKBUFX3 U439 ( .A(n15), .Y(n371) );
  CLKBUFX3 U440 ( .A(n501), .Y(n244) );
  CLKBUFX3 U441 ( .A(n509), .Y(n233) );
  CLKBUFX3 U442 ( .A(n509), .Y(n234) );
  CLKBUFX3 U443 ( .A(n206), .Y(n205) );
  CLKBUFX3 U444 ( .A(n365), .Y(n361) );
  CLKBUFX3 U445 ( .A(n501), .Y(n245) );
  CLKBUFX3 U446 ( .A(n11), .Y(n444) );
  CLKINVX1 U447 ( .A(n508), .Y(n238) );
  CLKINVX1 U448 ( .A(PCSrc), .Y(n1289) );
  CLKINVX1 U449 ( .A(n701), .Y(n1288) );
  AND4X1 U450 ( .A(n686), .B(ICACHE_rdata[27]), .C(n687), .D(n1288), .Y(n570)
         );
  NOR2X1 U451 ( .A(PCSrc), .B(ICACHE_rdata[28]), .Y(n687) );
  CLKBUFX3 U452 ( .A(n720), .Y(n229) );
  CLKBUFX3 U453 ( .A(n723), .Y(n222) );
  CLKBUFX3 U454 ( .A(n721), .Y(n227) );
  CLKBUFX3 U455 ( .A(n724), .Y(n219) );
  CLKBUFX3 U456 ( .A(n369), .Y(n353) );
  CLKBUFX3 U457 ( .A(n365), .Y(n363) );
  CLKBUFX3 U458 ( .A(n367), .Y(n357) );
  CLKBUFX3 U459 ( .A(n367), .Y(n359) );
  CLKINVX1 U460 ( .A(ICACHE_rdata[27]), .Y(n706) );
  CLKINVX1 U461 ( .A(ICACHE_rdata[28]), .Y(n705) );
  CLKBUFX3 U462 ( .A(n720), .Y(n230) );
  CLKBUFX3 U463 ( .A(n723), .Y(n224) );
  CLKBUFX3 U464 ( .A(n721), .Y(n228) );
  CLKBUFX3 U465 ( .A(n369), .Y(n355) );
  CLKBUFX3 U466 ( .A(n724), .Y(n220) );
  NOR3X1 U467 ( .A(ICACHE_rdata[30]), .B(ICACHE_rdata[31]), .C(
        ICACHE_rdata[29]), .Y(n686) );
  CLKINVX1 U468 ( .A(ICACHE_rdata[15]), .Y(n655) );
  CLKINVX1 U469 ( .A(ICACHE_rdata[14]), .Y(n656) );
  CLKINVX1 U470 ( .A(ICACHE_rdata[13]), .Y(n661) );
  CLKINVX1 U471 ( .A(ICACHE_rdata[12]), .Y(n662) );
  CLKINVX1 U472 ( .A(ICACHE_rdata[11]), .Y(n667) );
  CLKINVX1 U473 ( .A(ICACHE_rdata[10]), .Y(n668) );
  CLKINVX1 U474 ( .A(ICACHE_rdata[9]), .Y(n673) );
  CLKINVX1 U475 ( .A(ICACHE_rdata[8]), .Y(n674) );
  CLKINVX1 U476 ( .A(ICACHE_rdata[7]), .Y(n679) );
  CLKINVX1 U477 ( .A(ICACHE_rdata[6]), .Y(n680) );
  CLKINVX1 U478 ( .A(ICACHE_rdata[5]), .Y(n685) );
  CLKINVX1 U479 ( .A(ICACHE_rdata[4]), .Y(n688) );
  CLKINVX1 U480 ( .A(ICACHE_rdata[3]), .Y(n689) );
  CLKINVX1 U481 ( .A(ICACHE_rdata[2]), .Y(n694) );
  CLKINVX1 U482 ( .A(ICACHE_rdata[1]), .Y(n697) );
  CLKINVX1 U483 ( .A(ICACHE_rdata[0]), .Y(n698) );
  CLKBUFX3 U484 ( .A(n258), .Y(n279) );
  CLKBUFX3 U485 ( .A(n281), .Y(n285) );
  CLKBUFX3 U486 ( .A(n258), .Y(n281) );
  CLKBUFX3 U487 ( .A(n281), .Y(n283) );
  CLKBUFX3 U488 ( .A(n271), .Y(n273) );
  CLKBUFX3 U489 ( .A(n271), .Y(n277) );
  CLKBUFX3 U490 ( .A(n271), .Y(n275) );
  CLKBUFX3 U491 ( .A(n263), .Y(n265) );
  CLKBUFX3 U492 ( .A(n263), .Y(n269) );
  CLKBUFX3 U493 ( .A(n263), .Y(n267) );
  CLKINVX1 U494 ( .A(readreg2_forward[1]), .Y(n1530) );
  CLKBUFX3 U495 ( .A(n1534), .Y(n199) );
  CLKBUFX3 U496 ( .A(n1534), .Y(n200) );
  CLKINVX1 U497 ( .A(n456), .Y(n454) );
  CLKINVX1 U498 ( .A(readreg2_forward[0]), .Y(n1532) );
  CLKINVX1 U499 ( .A(readreg2_forward[5]), .Y(n1522) );
  CLKINVX1 U500 ( .A(readreg2_forward[4]), .Y(n1524) );
  CLKINVX1 U501 ( .A(readreg2_forward[8]), .Y(n1516) );
  CLKINVX1 U502 ( .A(readreg2_forward[7]), .Y(n1518) );
  CLKINVX1 U503 ( .A(readreg2_forward[6]), .Y(n1520) );
  CLKINVX1 U504 ( .A(readreg2_forward[3]), .Y(n1526) );
  CLKINVX1 U505 ( .A(readreg2_forward[2]), .Y(n1528) );
  CLKINVX1 U506 ( .A(readreg1_forward[4]), .Y(n1525) );
  CLKINVX1 U507 ( .A(readreg1_forward[3]), .Y(n1527) );
  CLKINVX1 U508 ( .A(readreg1_forward[2]), .Y(n1529) );
  CLKINVX1 U509 ( .A(readreg1_forward[0]), .Y(n1533) );
  CLKINVX1 U510 ( .A(readreg1_forward[1]), .Y(n1531) );
  OAI22XL U511 ( .A0(n203), .A1(n1548), .B0(n1524), .B1(n44), .Y(ALUin2[4]) );
  OAI22XL U512 ( .A0(n203), .A1(n1547), .B0(n1522), .B1(n206), .Y(ALUin2[5])
         );
  CLKBUFX3 U513 ( .A(n1535), .Y(n202) );
  CLKBUFX3 U514 ( .A(n1535), .Y(n201) );
  OAI22XL U515 ( .A0(n203), .A1(n1578), .B0(n1532), .B1(n207), .Y(ALUin2[0])
         );
  NOR3X1 U516 ( .A(stall_div), .B(stall_mul), .C(n319), .Y(n15) );
  NOR4X1 U517 ( .A(PCSrc), .B(ICACHE_rdata[27]), .C(n701), .D(n1470), .Y(n700)
         );
  CLKINVX1 U518 ( .A(readreg2_forward[16]), .Y(n1500) );
  CLKINVX1 U519 ( .A(readreg2_forward[15]), .Y(n1502) );
  CLKINVX1 U520 ( .A(readreg2_forward[14]), .Y(n1504) );
  CLKINVX1 U521 ( .A(readreg2_forward[13]), .Y(n1506) );
  CLKINVX1 U522 ( .A(readreg2_forward[12]), .Y(n1508) );
  CLKINVX1 U523 ( .A(readreg2_forward[11]), .Y(n1510) );
  CLKINVX1 U524 ( .A(readreg2_forward[10]), .Y(n1512) );
  CLKINVX1 U525 ( .A(readreg2_forward[9]), .Y(n1514) );
  NAND3X1 U526 ( .A(n708), .B(n1288), .C(n446), .Y(n13) );
  OAI21XL U527 ( .A0(n1550), .A1(n1538), .B0(IF_Flush), .Y(n708) );
  OA21X2 U528 ( .A0(n570), .A1(n571), .B0(n238), .Y(n550) );
  OAI22XL U529 ( .A0(n446), .A1(n1576), .B0(n437), .B1(n668), .Y(inst_w[10])
         );
  OAI22XL U530 ( .A0(n446), .A1(n1574), .B0(n439), .B1(n662), .Y(inst_w[12])
         );
  OAI22XL U531 ( .A0(n446), .A1(n1572), .B0(n441), .B1(n661), .Y(inst_w[13])
         );
  OAI22XL U532 ( .A0(n446), .A1(n1570), .B0(n439), .B1(n656), .Y(inst_w[14])
         );
  OAI22XL U533 ( .A0(n446), .A1(n45), .B0(n439), .B1(n655), .Y(inst_w[15]) );
  OAI22XL U534 ( .A0(n446), .A1(n1545), .B0(n437), .B1(n680), .Y(inst_w[6]) );
  OAI22XL U535 ( .A0(n446), .A1(n1543), .B0(n437), .B1(n679), .Y(inst_w[7]) );
  OAI22XL U536 ( .A0(n446), .A1(n1541), .B0(n437), .B1(n674), .Y(inst_w[8]) );
  OAI22XL U537 ( .A0(n446), .A1(n1539), .B0(n437), .B1(n673), .Y(inst_w[9]) );
  OAI22XL U538 ( .A0(n446), .A1(n1536), .B0(n439), .B1(n667), .Y(inst_w[11])
         );
  OAI22XL U539 ( .A0(n446), .A1(n1538), .B0(n437), .B1(n1470), .Y(take_w) );
  CLKBUFX3 U540 ( .A(n390), .Y(n252) );
  CLKBUFX3 U541 ( .A(n388), .Y(n256) );
  CLKBUFX3 U542 ( .A(n393), .Y(n250) );
  NAND3BX1 U543 ( .AN(stallJ), .B(PCWrite), .C(n387), .Y(n508) );
  CLKBUFX3 U544 ( .A(n393), .Y(n251) );
  CLKINVX1 U545 ( .A(n1389), .Y(n208) );
  CLKBUFX3 U546 ( .A(n388), .Y(n261) );
  NOR3BXL U547 ( .AN(IFIDWrite), .B(n389), .C(stallJ), .Y(n11) );
  NOR4BX1 U548 ( .AN(n693), .B(n1289), .C(n235), .D(JumpR), .Y(n503) );
  CLKINVX1 U549 ( .A(n295), .Y(n365) );
  NOR2BX1 U550 ( .AN(IF_Flush), .B(n1550), .Y(taken) );
  NOR3X1 U551 ( .A(n1550), .B(IF_Flush), .C(n1538), .Y(n701) );
  NAND2X1 U552 ( .A(raWrite), .B(n387), .Y(n498) );
  NOR4X1 U553 ( .A(n715), .B(n716), .C(n717), .D(n718), .Y(n714) );
  XOR2X1 U554 ( .A(n647), .B(n728), .Y(n715) );
  XOR2X1 U555 ( .A(n641), .B(n727), .Y(n716) );
  XOR2X1 U556 ( .A(n635), .B(n726), .Y(n717) );
  NOR4X1 U557 ( .A(n757), .B(n758), .C(n759), .D(n760), .Y(n756) );
  XOR2X1 U558 ( .A(n692), .B(n764), .Y(n757) );
  XOR2X1 U559 ( .A(n625), .B(n763), .Y(n758) );
  XOR2X1 U560 ( .A(n559), .B(n762), .Y(n759) );
  CLKINVX1 U561 ( .A(readreg2_forward[30]), .Y(n1472) );
  CLKINVX1 U562 ( .A(readreg2_forward[29]), .Y(n1474) );
  CLKINVX1 U563 ( .A(readreg2_forward[28]), .Y(n1476) );
  CLKINVX1 U564 ( .A(readreg2_forward[27]), .Y(n1478) );
  CLKINVX1 U565 ( .A(readreg2_forward[26]), .Y(n1480) );
  CLKINVX1 U566 ( .A(readreg2_forward[25]), .Y(n1482) );
  CLKINVX1 U567 ( .A(readreg2_forward[24]), .Y(n1484) );
  CLKINVX1 U568 ( .A(readreg2_forward[23]), .Y(n1486) );
  CLKINVX1 U569 ( .A(readreg2_forward[22]), .Y(n1488) );
  CLKINVX1 U570 ( .A(readreg2_forward[21]), .Y(n1490) );
  CLKINVX1 U571 ( .A(readreg2_forward[20]), .Y(n1492) );
  CLKINVX1 U572 ( .A(readreg2_forward[19]), .Y(n1494) );
  CLKINVX1 U573 ( .A(readreg2_forward[18]), .Y(n1496) );
  CLKINVX1 U574 ( .A(readreg2_forward[17]), .Y(n1498) );
  OAI22XL U575 ( .A0(n379), .A1(n1577), .B0(n410), .B1(n1576), .Y(
        sign_ext_w[10]) );
  OAI22XL U576 ( .A0(n379), .A1(n1546), .B0(n412), .B1(n1545), .Y(
        sign_ext_w[6]) );
  OAI22XL U577 ( .A0(n379), .A1(n1544), .B0(n412), .B1(n1543), .Y(
        sign_ext_w[7]) );
  OAI22XL U578 ( .A0(n375), .A1(n1542), .B0(n410), .B1(n1541), .Y(
        sign_ext_w[8]) );
  OAI22XL U579 ( .A0(n377), .A1(n1540), .B0(n398), .B1(n1539), .Y(
        sign_ext_w[9]) );
  OAI22XL U580 ( .A0(n379), .A1(n1575), .B0(n412), .B1(n1574), .Y(
        sign_ext_w[12]) );
  OAI22XL U581 ( .A0(n379), .A1(n1573), .B0(n412), .B1(n1572), .Y(
        sign_ext_w[13]) );
  OAI22XL U582 ( .A0(n381), .A1(n1571), .B0(n412), .B1(n1570), .Y(
        sign_ext_w[14]) );
  OAI22XL U583 ( .A0(n379), .A1(n1537), .B0(n410), .B1(n1536), .Y(
        sign_ext_w[11]) );
  OAI22XL U584 ( .A0(n377), .A1(n1643), .B0(n404), .B1(n1290), .Y(
        readreg1_w[31]) );
  OAI22XL U585 ( .A0(n377), .A1(n1642), .B0(n404), .B1(n1292), .Y(
        readreg1_w[30]) );
  OAI22XL U586 ( .A0(n377), .A1(n1641), .B0(n402), .B1(n1294), .Y(
        readreg1_w[29]) );
  OAI22XL U587 ( .A0(n381), .A1(n1640), .B0(n402), .B1(n1296), .Y(
        readreg1_w[28]) );
  OAI22XL U588 ( .A0(n383), .A1(n1639), .B0(n402), .B1(n1298), .Y(
        readreg1_w[27]) );
  OAI22XL U589 ( .A0(n375), .A1(n1638), .B0(n402), .B1(n1300), .Y(
        readreg1_w[26]) );
  OAI22XL U590 ( .A0(n381), .A1(n1637), .B0(n402), .B1(n1302), .Y(
        readreg1_w[25]) );
  OAI22XL U591 ( .A0(n383), .A1(n1636), .B0(n402), .B1(n1304), .Y(
        readreg1_w[24]) );
  OAI22XL U592 ( .A0(n375), .A1(n1635), .B0(n402), .B1(n1306), .Y(
        readreg1_w[23]) );
  OAI22XL U593 ( .A0(n379), .A1(n1634), .B0(n402), .B1(n1308), .Y(
        readreg1_w[22]) );
  OAI22XL U594 ( .A0(n377), .A1(n1633), .B0(n400), .B1(n1310), .Y(
        readreg1_w[21]) );
  OAI22XL U595 ( .A0(n381), .A1(n1632), .B0(n400), .B1(n1312), .Y(
        readreg1_w[20]) );
  OAI22XL U596 ( .A0(n383), .A1(n1631), .B0(n400), .B1(n1314), .Y(
        readreg1_w[19]) );
  OAI22XL U597 ( .A0(n375), .A1(n1630), .B0(n400), .B1(n1316), .Y(
        readreg1_w[18]) );
  OAI22XL U598 ( .A0(n379), .A1(n1629), .B0(n400), .B1(n1318), .Y(
        readreg1_w[17]) );
  OAI22XL U599 ( .A0(n375), .A1(n1628), .B0(n400), .B1(n1320), .Y(
        readreg1_w[16]) );
  OAI22XL U600 ( .A0(n375), .A1(n1627), .B0(n400), .B1(n1322), .Y(
        readreg1_w[15]) );
  OAI22XL U601 ( .A0(n375), .A1(n1626), .B0(n400), .B1(n1324), .Y(
        readreg1_w[14]) );
  OAI22XL U602 ( .A0(n375), .A1(n1625), .B0(n398), .B1(n1326), .Y(
        readreg1_w[13]) );
  OAI22XL U603 ( .A0(n375), .A1(n1624), .B0(n400), .B1(n1328), .Y(
        readreg1_w[12]) );
  OAI22XL U604 ( .A0(n375), .A1(n1623), .B0(n398), .B1(n1330), .Y(
        readreg1_w[11]) );
  OAI22XL U605 ( .A0(n375), .A1(n1622), .B0(n398), .B1(n1332), .Y(
        readreg1_w[10]) );
  OAI22XL U606 ( .A0(n377), .A1(n1621), .B0(n398), .B1(n1334), .Y(
        readreg1_w[9]) );
  OAI22XL U607 ( .A0(n377), .A1(n1620), .B0(n404), .B1(n1336), .Y(
        readreg1_w[8]) );
  OAI22XL U608 ( .A0(n377), .A1(n1619), .B0(n404), .B1(n1338), .Y(
        readreg1_w[7]) );
  OAI22XL U609 ( .A0(n377), .A1(n1618), .B0(n404), .B1(n1340), .Y(
        readreg1_w[6]) );
  OAI22XL U610 ( .A0(n377), .A1(n1617), .B0(n404), .B1(n1342), .Y(
        readreg1_w[5]) );
  OAI22XL U611 ( .A0(n377), .A1(n1616), .B0(n404), .B1(n1344), .Y(
        readreg1_w[4]) );
  OAI22XL U612 ( .A0(n377), .A1(n1615), .B0(n404), .B1(n1462), .Y(
        readreg1_w[3]) );
  OAI22XL U613 ( .A0(n377), .A1(n1614), .B0(n404), .B1(n1464), .Y(
        readreg1_w[2]) );
  OAI22XL U614 ( .A0(n377), .A1(n1613), .B0(n402), .B1(n1466), .Y(
        readreg1_w[1]) );
  OAI22XL U615 ( .A0(n375), .A1(n1612), .B0(n398), .B1(n1468), .Y(
        readreg1_w[0]) );
  OAI22XL U616 ( .A0(n381), .A1(n1611), .B0(n408), .B1(n1291), .Y(
        readreg2_w[31]) );
  OAI22XL U617 ( .A0(n381), .A1(n1610), .B0(n408), .B1(n1293), .Y(
        readreg2_w[30]) );
  OAI22XL U618 ( .A0(n381), .A1(n1609), .B0(n408), .B1(n1295), .Y(
        readreg2_w[29]) );
  OAI22XL U619 ( .A0(n381), .A1(n1608), .B0(n408), .B1(n1297), .Y(
        readreg2_w[28]) );
  OAI22XL U620 ( .A0(n381), .A1(n1607), .B0(n408), .B1(n1299), .Y(
        readreg2_w[27]) );
  OAI22XL U621 ( .A0(n383), .A1(n1606), .B0(n408), .B1(n1301), .Y(
        readreg2_w[26]) );
  OAI22XL U622 ( .A0(n383), .A1(n1605), .B0(n408), .B1(n1303), .Y(
        readreg2_w[25]) );
  OAI22XL U623 ( .A0(n383), .A1(n1604), .B0(n408), .B1(n1305), .Y(
        readreg2_w[24]) );
  OAI22XL U624 ( .A0(n383), .A1(n1603), .B0(n406), .B1(n1307), .Y(
        readreg2_w[23]) );
  OAI22XL U625 ( .A0(n383), .A1(n1602), .B0(n406), .B1(n1309), .Y(
        readreg2_w[22]) );
  OAI22XL U626 ( .A0(n383), .A1(n1601), .B0(n406), .B1(n1311), .Y(
        readreg2_w[21]) );
  OAI22XL U627 ( .A0(n383), .A1(n1600), .B0(n406), .B1(n1313), .Y(
        readreg2_w[20]) );
  OAI22XL U628 ( .A0(n383), .A1(n1599), .B0(n406), .B1(n1315), .Y(
        readreg2_w[19]) );
  OAI22XL U629 ( .A0(n383), .A1(n1598), .B0(n406), .B1(n1317), .Y(
        readreg2_w[18]) );
  OAI22XL U630 ( .A0(n375), .A1(n1597), .B0(n406), .B1(n1319), .Y(
        readreg2_w[17]) );
  OAI22XL U631 ( .A0(n383), .A1(n1596), .B0(n406), .B1(n1321), .Y(
        readreg2_w[16]) );
  OAI22XL U632 ( .A0(n379), .A1(n1595), .B0(n398), .B1(n1323), .Y(
        readreg2_w[15]) );
  OAI22XL U633 ( .A0(n377), .A1(n1594), .B0(n398), .B1(n1325), .Y(
        readreg2_w[14]) );
  OAI22XL U634 ( .A0(n383), .A1(n1593), .B0(n408), .B1(n1327), .Y(
        readreg2_w[13]) );
  OAI22XL U635 ( .A0(n383), .A1(n1592), .B0(n400), .B1(n1329), .Y(
        readreg2_w[12]) );
  OAI22XL U636 ( .A0(n381), .A1(n1591), .B0(n402), .B1(n1331), .Y(
        readreg2_w[11]) );
  OAI22XL U637 ( .A0(n383), .A1(n1590), .B0(n398), .B1(n1333), .Y(
        readreg2_w[10]) );
  OAI22XL U638 ( .A0(n379), .A1(n1589), .B0(n410), .B1(n1335), .Y(
        readreg2_w[9]) );
  OAI22XL U639 ( .A0(n381), .A1(n1588), .B0(n410), .B1(n1337), .Y(
        readreg2_w[8]) );
  OAI22XL U640 ( .A0(n381), .A1(n1587), .B0(n410), .B1(n1339), .Y(
        readreg2_w[7]) );
  OAI22XL U641 ( .A0(n381), .A1(n1586), .B0(n392), .B1(n1341), .Y(
        readreg2_w[6]) );
  OAI22XL U642 ( .A0(n381), .A1(n1585), .B0(n410), .B1(n1343), .Y(
        readreg2_w[5]) );
  OAI22XL U643 ( .A0(n381), .A1(n1584), .B0(n410), .B1(n1345), .Y(
        readreg2_w[4]) );
  OAI22XL U644 ( .A0(n381), .A1(n1583), .B0(n410), .B1(n1463), .Y(
        readreg2_w[3]) );
  OAI22XL U645 ( .A0(n381), .A1(n1582), .B0(n408), .B1(n1465), .Y(
        readreg2_w[2]) );
  OAI22XL U646 ( .A0(n383), .A1(n1581), .B0(n406), .B1(n1467), .Y(
        readreg2_w[1]) );
  OAI22XL U647 ( .A0(n377), .A1(n1580), .B0(n408), .B1(n1469), .Y(
        readreg2_w[0]) );
  NAND4X1 U648 ( .A(n711), .B(n712), .C(n713), .D(n714), .Y(n710) );
  NOR4X1 U649 ( .A(n737), .B(n738), .C(n739), .D(n740), .Y(n712) );
  NOR4X1 U650 ( .A(n729), .B(n730), .C(n731), .D(n732), .Y(n713) );
  NOR4X1 U651 ( .A(n745), .B(n746), .C(n747), .D(n748), .Y(n711) );
  NAND4X1 U652 ( .A(n753), .B(n754), .C(n755), .D(n756), .Y(n709) );
  NOR4X1 U653 ( .A(n781), .B(n782), .C(n783), .D(n784), .Y(n753) );
  NOR4X1 U654 ( .A(n773), .B(n774), .C(n775), .D(n776), .Y(n754) );
  NOR4X1 U655 ( .A(n765), .B(n766), .C(n767), .D(n768), .Y(n755) );
  CLKINVX1 U656 ( .A(PC_4[27]), .Y(n572) );
  CLKINVX1 U657 ( .A(PC_4[26]), .Y(n573) );
  CLKBUFX3 U658 ( .A(n29), .Y(n197) );
  NAND2X1 U659 ( .A(n198), .B(n387), .Y(n29) );
  OAI2BB2XL U660 ( .B0(n373), .B1(n203), .A0N(ALUSrc), .A1N(n196), .Y(
        ALUSrc_idex_w) );
  OAI21XL U661 ( .A0(n373), .A1(n1567), .B0(n197), .Y(sign_ext_w[17]) );
  OAI21XL U662 ( .A0(n373), .A1(n1565), .B0(n197), .Y(sign_ext_w[19]) );
  OAI21XL U663 ( .A0(n373), .A1(n1564), .B0(n197), .Y(sign_ext_w[20]) );
  OAI21XL U664 ( .A0(n373), .A1(n1563), .B0(n197), .Y(sign_ext_w[21]) );
  OAI21XL U665 ( .A0(n373), .A1(n1562), .B0(n197), .Y(sign_ext_w[22]) );
  OAI21XL U666 ( .A0(n373), .A1(n1561), .B0(n197), .Y(sign_ext_w[23]) );
  OAI21XL U667 ( .A0(n373), .A1(n1560), .B0(n197), .Y(sign_ext_w[24]) );
  OAI21XL U668 ( .A0(n373), .A1(n1558), .B0(n197), .Y(sign_ext_w[26]) );
  OAI21XL U669 ( .A0(n373), .A1(n1557), .B0(n197), .Y(sign_ext_w[27]) );
  OAI21XL U670 ( .A0(n373), .A1(n1556), .B0(n197), .Y(sign_ext_w[28]) );
  OAI21XL U671 ( .A0(n373), .A1(n1555), .B0(n197), .Y(sign_ext_w[29]) );
  OAI21XL U672 ( .A0(n373), .A1(n1554), .B0(n197), .Y(sign_ext_w[30]) );
  OAI21XL U673 ( .A0(n373), .A1(n1553), .B0(n197), .Y(sign_ext_w[31]) );
  OAI21XL U674 ( .A0(n375), .A1(n1569), .B0(n197), .Y(sign_ext_w[15]) );
  OAI21XL U675 ( .A0(n375), .A1(n1568), .B0(n197), .Y(sign_ext_w[16]) );
  OAI21XL U676 ( .A0(n375), .A1(n1566), .B0(n197), .Y(sign_ext_w[18]) );
  OAI21XL U677 ( .A0(n375), .A1(n1559), .B0(n197), .Y(sign_ext_w[25]) );
  CLKINVX1 U678 ( .A(Readdata1[30]), .Y(n1292) );
  CLKINVX1 U679 ( .A(Readdata1[9]), .Y(n1334) );
  CLKINVX1 U680 ( .A(Readdata1[7]), .Y(n1338) );
  CLKINVX1 U681 ( .A(Readdata1[6]), .Y(n1340) );
  CLKINVX1 U682 ( .A(Readdata1[5]), .Y(n1342) );
  CLKINVX1 U683 ( .A(Readdata1[3]), .Y(n1462) );
  CLKINVX1 U684 ( .A(Readdata2[19]), .Y(n1315) );
  CLKINVX1 U685 ( .A(Readdata1[31]), .Y(n1290) );
  CLKINVX1 U686 ( .A(Readdata1[29]), .Y(n1294) );
  CLKINVX1 U687 ( .A(Readdata1[27]), .Y(n1298) );
  CLKINVX1 U688 ( .A(Readdata1[26]), .Y(n1300) );
  CLKINVX1 U689 ( .A(Readdata1[25]), .Y(n1302) );
  CLKINVX1 U690 ( .A(Readdata1[23]), .Y(n1306) );
  CLKINVX1 U691 ( .A(Readdata1[22]), .Y(n1308) );
  CLKINVX1 U692 ( .A(Readdata1[21]), .Y(n1310) );
  CLKINVX1 U693 ( .A(Readdata1[19]), .Y(n1314) );
  CLKINVX1 U694 ( .A(Readdata1[18]), .Y(n1316) );
  CLKINVX1 U695 ( .A(Readdata1[17]), .Y(n1318) );
  CLKINVX1 U696 ( .A(Readdata1[15]), .Y(n1322) );
  CLKINVX1 U697 ( .A(Readdata1[14]), .Y(n1324) );
  CLKINVX1 U698 ( .A(Readdata1[13]), .Y(n1326) );
  CLKINVX1 U699 ( .A(Readdata1[11]), .Y(n1330) );
  CLKINVX1 U700 ( .A(Readdata1[10]), .Y(n1332) );
  CLKINVX1 U701 ( .A(Readdata1[2]), .Y(n1464) );
  CLKINVX1 U702 ( .A(Readdata1[1]), .Y(n1466) );
  CLKINVX1 U703 ( .A(Readdata1[0]), .Y(n1468) );
  CLKBUFX3 U704 ( .A(n390), .Y(n255) );
  CLKBUFX3 U705 ( .A(n223), .Y(n287) );
  CLKBUFX3 U706 ( .A(n223), .Y(n289) );
  CLKBUFX3 U707 ( .A(n497), .Y(n196) );
  NOR3X1 U708 ( .A(stall), .B(stallJ), .C(n397), .Y(n497) );
  CLKBUFX3 U709 ( .A(n221), .Y(n293) );
  CLKBUFX3 U710 ( .A(n221), .Y(n291) );
  CLKINVX1 U711 ( .A(n295), .Y(n367) );
  CLKINVX1 U712 ( .A(n295), .Y(n369) );
  CLKINVX1 U713 ( .A(n396), .Y(n1461) );
  CLKINVX1 U714 ( .A(n450), .Y(n1458) );
  CLKINVX1 U715 ( .A(n453), .Y(n1457) );
  CLKINVX1 U716 ( .A(n455), .Y(n1456) );
  CLKINVX1 U717 ( .A(n457), .Y(n1455) );
  CLKINVX1 U718 ( .A(n459), .Y(n1454) );
  CLKINVX1 U719 ( .A(n461), .Y(n1453) );
  CLKINVX1 U720 ( .A(n463), .Y(n1452) );
  CLKINVX1 U721 ( .A(n399), .Y(n1451) );
  CLKINVX1 U722 ( .A(n401), .Y(n1450) );
  CLKINVX1 U723 ( .A(n415), .Y(n1443) );
  CLKINVX1 U724 ( .A(n447), .Y(n1430) );
  CLKINVX1 U725 ( .A(PC_4[25]), .Y(n578) );
  CLKINVX1 U726 ( .A(PC_4[24]), .Y(n579) );
  CLKINVX1 U727 ( .A(PC_4[23]), .Y(n584) );
  CLKINVX1 U728 ( .A(PC_4[22]), .Y(n585) );
  CLKINVX1 U729 ( .A(PC_4[21]), .Y(n590) );
  CLKINVX1 U730 ( .A(PC_4[20]), .Y(n591) );
  CLKINVX1 U731 ( .A(PC_4[19]), .Y(n596) );
  CLKINVX1 U732 ( .A(PC_4[18]), .Y(n597) );
  CLKINVX1 U733 ( .A(n420), .Y(n1460) );
  CLKINVX1 U734 ( .A(n443), .Y(n1459) );
  CLKINVX1 U735 ( .A(n403), .Y(n1449) );
  CLKINVX1 U736 ( .A(n405), .Y(n1448) );
  CLKINVX1 U737 ( .A(n407), .Y(n1447) );
  CLKINVX1 U738 ( .A(n409), .Y(n1446) );
  CLKINVX1 U739 ( .A(n411), .Y(n1445) );
  CLKINVX1 U740 ( .A(n413), .Y(n1444) );
  CLKINVX1 U741 ( .A(n417), .Y(n1442) );
  CLKINVX1 U742 ( .A(n422), .Y(n1441) );
  CLKINVX1 U743 ( .A(n424), .Y(n1440) );
  CLKINVX1 U744 ( .A(n426), .Y(n1439) );
  CLKINVX1 U745 ( .A(n428), .Y(n1438) );
  CLKINVX1 U746 ( .A(n430), .Y(n1437) );
  CLKINVX1 U747 ( .A(n432), .Y(n1436) );
  CLKINVX1 U748 ( .A(n434), .Y(n1435) );
  CLKINVX1 U749 ( .A(n436), .Y(n1434) );
  CLKINVX1 U750 ( .A(n438), .Y(n1433) );
  CLKINVX1 U751 ( .A(n440), .Y(n1432) );
  CLKINVX1 U752 ( .A(n445), .Y(n1431) );
  CLKINVX1 U753 ( .A(Readdata2[30]), .Y(n1293) );
  CLKINVX1 U754 ( .A(Readdata2[3]), .Y(n1463) );
  CLKINVX1 U755 ( .A(Readdata2[7]), .Y(n1339) );
  CLKINVX1 U756 ( .A(Readdata2[6]), .Y(n1341) );
  CLKINVX1 U757 ( .A(Readdata2[5]), .Y(n1343) );
  CLKINVX1 U758 ( .A(Readdata2[4]), .Y(n1345) );
  CLKINVX1 U759 ( .A(Readdata2[9]), .Y(n1335) );
  CLKINVX1 U760 ( .A(Readdata2[8]), .Y(n1337) );
  CLKINVX1 U761 ( .A(Readdata1[8]), .Y(n1336) );
  CLKINVX1 U762 ( .A(Readdata1[4]), .Y(n1344) );
  CLKINVX1 U763 ( .A(Readdata2[18]), .Y(n1317) );
  CLKINVX1 U764 ( .A(Readdata2[17]), .Y(n1319) );
  CLKINVX1 U765 ( .A(Readdata2[16]), .Y(n1321) );
  CLKINVX1 U766 ( .A(Readdata2[31]), .Y(n1291) );
  CLKINVX1 U767 ( .A(Readdata2[29]), .Y(n1295) );
  CLKINVX1 U768 ( .A(Readdata1[28]), .Y(n1296) );
  CLKINVX1 U769 ( .A(Readdata2[28]), .Y(n1297) );
  CLKINVX1 U770 ( .A(Readdata2[23]), .Y(n1307) );
  CLKINVX1 U771 ( .A(Readdata2[22]), .Y(n1309) );
  CLKINVX1 U772 ( .A(Readdata2[21]), .Y(n1311) );
  CLKINVX1 U773 ( .A(Readdata2[20]), .Y(n1313) );
  CLKINVX1 U774 ( .A(Readdata2[26]), .Y(n1301) );
  CLKINVX1 U775 ( .A(Readdata2[27]), .Y(n1299) );
  CLKINVX1 U776 ( .A(Readdata2[25]), .Y(n1303) );
  CLKINVX1 U777 ( .A(Readdata2[24]), .Y(n1305) );
  CLKINVX1 U778 ( .A(Readdata2[2]), .Y(n1465) );
  CLKINVX1 U779 ( .A(Readdata2[1]), .Y(n1467) );
  CLKINVX1 U780 ( .A(Readdata2[11]), .Y(n1331) );
  CLKINVX1 U781 ( .A(Readdata2[10]), .Y(n1333) );
  CLKINVX1 U782 ( .A(Readdata2[15]), .Y(n1323) );
  CLKINVX1 U783 ( .A(Readdata2[14]), .Y(n1325) );
  CLKINVX1 U784 ( .A(Readdata2[13]), .Y(n1327) );
  CLKINVX1 U785 ( .A(Readdata2[12]), .Y(n1329) );
  CLKINVX1 U786 ( .A(Readdata1[24]), .Y(n1304) );
  CLKINVX1 U787 ( .A(Readdata1[20]), .Y(n1312) );
  CLKINVX1 U788 ( .A(Readdata1[16]), .Y(n1320) );
  CLKINVX1 U789 ( .A(Readdata1[12]), .Y(n1328) );
  CLKINVX1 U790 ( .A(Readdata2[0]), .Y(n1469) );
  CLKINVX1 U791 ( .A(Branch), .Y(n1550) );
  CLKINVX1 U792 ( .A(ICACHE_rdata[25]), .Y(n789) );
  CLKINVX1 U793 ( .A(ICACHE_rdata[24]), .Y(n791) );
  CLKINVX1 U794 ( .A(ICACHE_rdata[23]), .Y(n915) );
  CLKINVX1 U795 ( .A(ICACHE_rdata[22]), .Y(n916) );
  CLKINVX1 U796 ( .A(ICACHE_rdata[21]), .Y(n917) );
  CLKINVX1 U797 ( .A(ICACHE_rdata[20]), .Y(n918) );
  CLKINVX1 U798 ( .A(ICACHE_rdata[19]), .Y(n919) );
  CLKINVX1 U799 ( .A(ICACHE_rdata[18]), .Y(n920) );
  CLKINVX1 U800 ( .A(ICACHE_rdata[17]), .Y(n649) );
  CLKINVX1 U801 ( .A(ICACHE_rdata[16]), .Y(n650) );
  CLKINVX1 U802 ( .A(PC_4[17]), .Y(n602) );
  CLKINVX1 U803 ( .A(PC_4[16]), .Y(n603) );
  CLKINVX1 U804 ( .A(PC_4[15]), .Y(n608) );
  CLKINVX1 U805 ( .A(PC_4[14]), .Y(n609) );
  CLKINVX1 U806 ( .A(PC_4[13]), .Y(n614) );
  CLKINVX1 U807 ( .A(PC_4[12]), .Y(n615) );
  CLKINVX1 U808 ( .A(PC_4[11]), .Y(n620) );
  CLKINVX1 U809 ( .A(PC_4[10]), .Y(n621) );
  CLKINVX1 U810 ( .A(PC_4[3]), .Y(n643) );
  CLKINVX1 U811 ( .A(PC_4[6]), .Y(n632) );
  CLKINVX1 U812 ( .A(PC_4[5]), .Y(n637) );
  CLKINVX1 U813 ( .A(PC_4[4]), .Y(n638) );
  CLKINVX1 U814 ( .A(PC_4[9]), .Y(n624) );
  CLKINVX1 U815 ( .A(PC_4[8]), .Y(n626) );
  CLKINVX1 U816 ( .A(PC_4[7]), .Y(n631) );
  OAI222XL U817 ( .A0(n309), .A1(n1398), .B0(n291), .B1(n1103), .C0(n481), 
        .C1(n287), .Y(n1248) );
  CLKINVX1 U818 ( .A(ALUresult[31]), .Y(n481) );
  OAI222XL U819 ( .A0(n1611), .A1(n215), .B0(n200), .B1(n447), .C0(n1398), 
        .C1(n213), .Y(readreg2_forward[31]) );
  OAI222XL U820 ( .A0(n311), .A1(n1399), .B0(n291), .B1(n1018), .C0(n482), 
        .C1(n287), .Y(n1171) );
  CLKINVX1 U821 ( .A(ALUresult[30]), .Y(n482) );
  OAI222XL U822 ( .A0(n313), .A1(n1401), .B0(n293), .B1(n1022), .C0(n484), 
        .C1(n287), .Y(n1175) );
  CLKINVX1 U823 ( .A(ALUresult[28]), .Y(n484) );
  OAI222XL U824 ( .A0(n313), .A1(n1403), .B0(n221), .B1(n1026), .C0(n486), 
        .C1(n287), .Y(n1179) );
  CLKINVX1 U825 ( .A(ALUresult[26]), .Y(n486) );
  OAI222XL U826 ( .A0(n311), .A1(n1405), .B0(n221), .B1(n1030), .C0(n488), 
        .C1(n287), .Y(n1183) );
  CLKINVX1 U827 ( .A(ALUresult[24]), .Y(n488) );
  OAI222XL U828 ( .A0(n309), .A1(n1402), .B0(n221), .B1(n1024), .C0(n485), 
        .C1(n287), .Y(n1177) );
  CLKINVX1 U829 ( .A(ALUresult[27]), .Y(n485) );
  OAI222XL U830 ( .A0(n311), .A1(n1404), .B0(n221), .B1(n1028), .C0(n487), 
        .C1(n287), .Y(n1181) );
  CLKINVX1 U831 ( .A(ALUresult[25]), .Y(n487) );
  OAI222XL U832 ( .A0(n311), .A1(n1400), .B0(n291), .B1(n1020), .C0(n483), 
        .C1(n287), .Y(n1173) );
  CLKINVX1 U833 ( .A(ALUresult[29]), .Y(n483) );
  CLKBUFX3 U834 ( .A(n1105), .Y(n211) );
  CLKBUFX3 U835 ( .A(n1105), .Y(n209) );
  CLKBUFX3 U836 ( .A(n1105), .Y(n210) );
  OAI222XL U837 ( .A0(n1521), .A1(n252), .B0(n828), .B1(n261), .C0(n861), .C1(
        n250), .Y(n1374) );
  CLKINVX1 U838 ( .A(readreg1_forward[6]), .Y(n1521) );
  OAI222XL U839 ( .A0(n1523), .A1(n252), .B0(n827), .B1(n261), .C0(n860), .C1(
        n250), .Y(n1373) );
  CLKINVX1 U840 ( .A(readreg1_forward[5]), .Y(n1523) );
  OAI222XL U841 ( .A0(n311), .A1(n1406), .B0(n293), .B1(n1032), .C0(n489), 
        .C1(n287), .Y(n1185) );
  CLKINVX1 U842 ( .A(ALUresult[23]), .Y(n489) );
  OAI221XL U843 ( .A0(n800), .A1(n256), .B0(n1533), .B1(n252), .C0(n391), .Y(
        n1346) );
  AOI2BB2X1 U844 ( .B0(shamt_idex_r[0]), .B1(n43), .A0N(n833), .A1N(n251), .Y(
        n391) );
  OAI221XL U845 ( .A0(n826), .A1(n256), .B0(n1525), .B1(n252), .C0(n452), .Y(
        n1372) );
  AOI2BB2X1 U846 ( .B0(shamt_idex_r[4]), .B1(n43), .A0N(n859), .A1N(n251), .Y(
        n452) );
  OAI221XL U847 ( .A0(n825), .A1(n256), .B0(n1527), .B1(n252), .C0(n449), .Y(
        n1371) );
  AOI2BB2X1 U848 ( .B0(shamt_idex_r[3]), .B1(n43), .A0N(n858), .A1N(n251), .Y(
        n449) );
  OAI221XL U849 ( .A0(n822), .A1(n256), .B0(n1529), .B1(n252), .C0(n442), .Y(
        n1368) );
  AOI2BB2X1 U850 ( .B0(shamt_idex_r[2]), .B1(n43), .A0N(n855), .A1N(n251), .Y(
        n442) );
  OAI221XL U851 ( .A0(n811), .A1(n256), .B0(n1531), .B1(n252), .C0(n419), .Y(
        n1357) );
  AOI2BB2X1 U852 ( .B0(shamt_idex_r[1]), .B1(n43), .A0N(n844), .A1N(n251), .Y(
        n419) );
  OAI222XL U853 ( .A0(n311), .A1(n1407), .B0(n293), .B1(n1034), .C0(n490), 
        .C1(n287), .Y(n1187) );
  CLKINVX1 U854 ( .A(ALUresult[22]), .Y(n490) );
  OAI222XL U855 ( .A0(n311), .A1(n1409), .B0(n293), .B1(n1038), .C0(n492), 
        .C1(n287), .Y(n1191) );
  CLKINVX1 U856 ( .A(ALUresult[20]), .Y(n492) );
  OAI222XL U857 ( .A0(n311), .A1(n1410), .B0(n293), .B1(n1040), .C0(n493), 
        .C1(n287), .Y(n1193) );
  CLKINVX1 U858 ( .A(ALUresult[19]), .Y(n493) );
  OAI222XL U859 ( .A0(n311), .A1(n1412), .B0(n293), .B1(n1044), .C0(n495), 
        .C1(n289), .Y(n1197) );
  CLKINVX1 U860 ( .A(ALUresult[17]), .Y(n495) );
  OAI222XL U861 ( .A0(n311), .A1(n1413), .B0(n293), .B1(n1046), .C0(n496), 
        .C1(n289), .Y(n1199) );
  CLKINVX1 U862 ( .A(ALUresult[16]), .Y(n496) );
  NAND2X1 U863 ( .A(n574), .B(n575), .Y(PC_w[27]) );
  AOI222XL U864 ( .A0(n236), .A1(ICACHE_addr[25]), .B0(N113), .B1(n234), .C0(
        n232), .C1(PC_4_r[27]), .Y(n574) );
  AOI221XL U865 ( .A0(n244), .A1(n576), .B0(N325), .B1(n243), .C0(n577), .Y(
        n575) );
  NAND2X1 U866 ( .A(n580), .B(n581), .Y(PC_w[26]) );
  AOI222XL U867 ( .A0(n236), .A1(ICACHE_addr[24]), .B0(N112), .B1(n234), .C0(
        n232), .C1(PC_4_r[26]), .Y(n580) );
  AOI221XL U868 ( .A0(n244), .A1(n582), .B0(N324), .B1(n243), .C0(n583), .Y(
        n581) );
  NAND2X1 U869 ( .A(n586), .B(n587), .Y(PC_w[25]) );
  AOI222XL U870 ( .A0(n236), .A1(ICACHE_addr[23]), .B0(N111), .B1(n234), .C0(
        n232), .C1(PC_4_r[25]), .Y(n586) );
  AOI221XL U871 ( .A0(n244), .A1(n588), .B0(N323), .B1(n243), .C0(n589), .Y(
        n587) );
  NAND2X1 U872 ( .A(n592), .B(n593), .Y(PC_w[24]) );
  AOI222XL U873 ( .A0(n236), .A1(ICACHE_addr[22]), .B0(N110), .B1(n234), .C0(
        n232), .C1(PC_4_r[24]), .Y(n592) );
  AOI221XL U874 ( .A0(n244), .A1(n594), .B0(N322), .B1(n243), .C0(n595), .Y(
        n593) );
  NAND2X1 U875 ( .A(n598), .B(n599), .Y(PC_w[23]) );
  AOI222XL U876 ( .A0(n236), .A1(ICACHE_addr[21]), .B0(N109), .B1(n234), .C0(
        n232), .C1(PC_4_r[23]), .Y(n598) );
  AOI221XL U877 ( .A0(n244), .A1(n600), .B0(N321), .B1(n243), .C0(n601), .Y(
        n599) );
  NAND2X1 U878 ( .A(n604), .B(n605), .Y(PC_w[22]) );
  AOI222XL U879 ( .A0(n236), .A1(ICACHE_addr[20]), .B0(N108), .B1(n233), .C0(
        n232), .C1(PC_4_r[22]), .Y(n604) );
  AOI221XL U880 ( .A0(n244), .A1(n606), .B0(N320), .B1(n243), .C0(n607), .Y(
        n605) );
  NAND2X1 U881 ( .A(n610), .B(n611), .Y(PC_w[21]) );
  AOI222XL U882 ( .A0(n235), .A1(ICACHE_addr[19]), .B0(N107), .B1(n234), .C0(
        n232), .C1(PC_4_r[21]), .Y(n610) );
  AOI221XL U883 ( .A0(n244), .A1(n612), .B0(N319), .B1(n243), .C0(n613), .Y(
        n611) );
  NAND2X1 U884 ( .A(n616), .B(n617), .Y(PC_w[20]) );
  AOI222XL U885 ( .A0(n235), .A1(ICACHE_addr[18]), .B0(N106), .B1(n233), .C0(
        n232), .C1(PC_4_r[20]), .Y(n616) );
  AOI221XL U886 ( .A0(n244), .A1(n618), .B0(N318), .B1(n243), .C0(n619), .Y(
        n617) );
  NAND2X1 U887 ( .A(n627), .B(n628), .Y(PC_w[19]) );
  AOI222XL U888 ( .A0(n235), .A1(ICACHE_addr[17]), .B0(N105), .B1(n234), .C0(
        n232), .C1(PC_4_r[19]), .Y(n627) );
  AOI221XL U889 ( .A0(n244), .A1(n629), .B0(N317), .B1(n243), .C0(n630), .Y(
        n628) );
  NAND2X1 U890 ( .A(n633), .B(n634), .Y(PC_w[18]) );
  AOI222XL U891 ( .A0(n235), .A1(ICACHE_addr[16]), .B0(N104), .B1(n233), .C0(
        n232), .C1(PC_4_r[18]), .Y(n633) );
  AOI221XL U892 ( .A0(n244), .A1(n635), .B0(N316), .B1(n243), .C0(n636), .Y(
        n634) );
  NAND2X1 U893 ( .A(n639), .B(n640), .Y(PC_w[17]) );
  AOI222XL U894 ( .A0(n235), .A1(ICACHE_addr[15]), .B0(N103), .B1(n509), .C0(
        n232), .C1(PC_4_r[17]), .Y(n639) );
  AOI221XL U895 ( .A0(n244), .A1(n641), .B0(N315), .B1(n243), .C0(n642), .Y(
        n640) );
  NAND2X1 U896 ( .A(n657), .B(n658), .Y(PC_w[14]) );
  AOI222XL U897 ( .A0(n235), .A1(ICACHE_addr[12]), .B0(N100), .B1(n234), .C0(
        n232), .C1(PC_4_r[14]), .Y(n657) );
  AOI221XL U898 ( .A0(n244), .A1(n659), .B0(N312), .B1(n243), .C0(n660), .Y(
        n658) );
  NAND2X1 U899 ( .A(n557), .B(n558), .Y(PC_w[2]) );
  AOI222XL U900 ( .A0(n236), .A1(ICACHE_addr[0]), .B0(N88), .B1(n233), .C0(
        n231), .C1(PC_4_r[2]), .Y(n557) );
  AOI221XL U901 ( .A0(n244), .A1(n559), .B0(N300), .B1(n243), .C0(n560), .Y(
        n558) );
  OAI22XL U902 ( .A0(n240), .A1(ICACHE_addr[0]), .B0(n698), .B1(n239), .Y(n560) );
  OAI22XL U903 ( .A0(n890), .A1(n448), .B0(n439), .B1(ICACHE_addr[0]), .Y(
        PC_4_w[2]) );
  OAI22XL U904 ( .A0(n910), .A1(n451), .B0(n441), .B1(n706), .Y(inst_w[27]) );
  OAI22XL U905 ( .A0(n911), .A1(n451), .B0(n441), .B1(n705), .Y(inst_w[28]) );
  OAI22XL U906 ( .A0(n948), .A1(n451), .B0(n441), .B1(n697), .Y(inst_w[1]) );
  OAI22XL U907 ( .A0(n949), .A1(n451), .B0(n441), .B1(n694), .Y(inst_w[2]) );
  OAI22XL U908 ( .A0(n950), .A1(n451), .B0(n441), .B1(n689), .Y(inst_w[3]) );
  OAI22XL U909 ( .A0(n951), .A1(n448), .B0(n441), .B1(n688), .Y(inst_w[4]) );
  OAI22XL U910 ( .A0(n952), .A1(n448), .B0(n441), .B1(n685), .Y(inst_w[5]) );
  OAI22XL U911 ( .A0(n947), .A1(n451), .B0(n441), .B1(n698), .Y(inst_w[0]) );
  OAI22XL U912 ( .A0(n1388), .A1(n451), .B0(n441), .B1(n650), .Y(inst_w[16])
         );
  OAI22XL U913 ( .A0(n1387), .A1(n451), .B0(n439), .B1(n649), .Y(inst_w[17])
         );
  OAI22XL U914 ( .A0(n1386), .A1(n451), .B0(n441), .B1(n920), .Y(inst_w[18])
         );
  OAI22XL U915 ( .A0(n1385), .A1(n451), .B0(n439), .B1(n919), .Y(inst_w[19])
         );
  OAI22XL U916 ( .A0(n1384), .A1(n451), .B0(n439), .B1(n918), .Y(inst_w[20])
         );
  OAI22XL U917 ( .A0(n904), .A1(n451), .B0(n441), .B1(n917), .Y(inst_w[21]) );
  OAI22XL U918 ( .A0(n905), .A1(n451), .B0(n441), .B1(n916), .Y(inst_w[22]) );
  OAI22XL U919 ( .A0(n906), .A1(n451), .B0(n441), .B1(n915), .Y(inst_w[23]) );
  OAI22XL U920 ( .A0(n907), .A1(n451), .B0(n441), .B1(n791), .Y(inst_w[24]) );
  OAI22XL U921 ( .A0(n908), .A1(n451), .B0(n441), .B1(n789), .Y(inst_w[25]) );
  OAI22XL U922 ( .A0(n889), .A1(n451), .B0(n439), .B1(n572), .Y(PC_4_w[27]) );
  OAI22XL U923 ( .A0(n888), .A1(n448), .B0(n439), .B1(n573), .Y(PC_4_w[26]) );
  OAI22XL U924 ( .A0(n887), .A1(n451), .B0(n439), .B1(n578), .Y(PC_4_w[25]) );
  OAI22XL U925 ( .A0(n886), .A1(n448), .B0(n439), .B1(n579), .Y(PC_4_w[24]) );
  OAI22XL U926 ( .A0(n885), .A1(n451), .B0(n439), .B1(n584), .Y(PC_4_w[23]) );
  OAI22XL U927 ( .A0(n884), .A1(n448), .B0(n439), .B1(n585), .Y(PC_4_w[22]) );
  OAI22XL U928 ( .A0(n883), .A1(n448), .B0(n439), .B1(n590), .Y(PC_4_w[21]) );
  OAI22XL U929 ( .A0(n882), .A1(n448), .B0(n439), .B1(n591), .Y(PC_4_w[20]) );
  OAI22XL U930 ( .A0(n881), .A1(n448), .B0(n437), .B1(n596), .Y(PC_4_w[19]) );
  OAI22XL U931 ( .A0(n880), .A1(n448), .B0(n437), .B1(n597), .Y(PC_4_w[18]) );
  OAI22XL U932 ( .A0(n891), .A1(n451), .B0(n437), .B1(n643), .Y(PC_4_w[3]) );
  OAI22XL U933 ( .A0(n914), .A1(n448), .B0(n441), .B1(n699), .Y(inst_w[31]) );
  CLKINVX1 U934 ( .A(ICACHE_rdata[31]), .Y(n699) );
  OAI22XL U935 ( .A0(n912), .A1(n448), .B0(n441), .B1(n704), .Y(inst_w[29]) );
  CLKINVX1 U936 ( .A(ICACHE_rdata[29]), .Y(n704) );
  OAI22XL U937 ( .A0(n913), .A1(n448), .B0(n441), .B1(n703), .Y(inst_w[30]) );
  CLKINVX1 U938 ( .A(ICACHE_rdata[30]), .Y(n703) );
  OAI22XL U939 ( .A0(n879), .A1(n448), .B0(n437), .B1(n602), .Y(PC_4_w[17]) );
  OAI22XL U940 ( .A0(n878), .A1(n448), .B0(n437), .B1(n603), .Y(PC_4_w[16]) );
  OAI22XL U941 ( .A0(n877), .A1(n448), .B0(n437), .B1(n608), .Y(PC_4_w[15]) );
  OAI22XL U942 ( .A0(n876), .A1(n446), .B0(n437), .B1(n609), .Y(PC_4_w[14]) );
  OAI22XL U943 ( .A0(n875), .A1(n448), .B0(n437), .B1(n614), .Y(PC_4_w[13]) );
  OAI22XL U944 ( .A0(n874), .A1(n448), .B0(n437), .B1(n615), .Y(PC_4_w[12]) );
  OAI22XL U945 ( .A0(n873), .A1(n446), .B0(n437), .B1(n620), .Y(PC_4_w[11]) );
  OAI22XL U946 ( .A0(n872), .A1(n448), .B0(n437), .B1(n621), .Y(PC_4_w[10]) );
  OAI22XL U947 ( .A0(n897), .A1(n446), .B0(n13), .B1(n624), .Y(PC_4_w[9]) );
  OAI22XL U948 ( .A0(n896), .A1(n444), .B0(n13), .B1(n626), .Y(PC_4_w[8]) );
  OAI22XL U949 ( .A0(n895), .A1(n444), .B0(n13), .B1(n631), .Y(PC_4_w[7]) );
  OAI22XL U950 ( .A0(n894), .A1(n444), .B0(n439), .B1(n632), .Y(PC_4_w[6]) );
  OAI22XL U951 ( .A0(n893), .A1(n444), .B0(n441), .B1(n637), .Y(PC_4_w[5]) );
  OAI22XL U952 ( .A0(n892), .A1(n444), .B0(n437), .B1(n638), .Y(PC_4_w[4]) );
  OAI22XL U953 ( .A0(n1379), .A1(n444), .B0(n439), .B1(n561), .Y(PC_4_w[30])
         );
  CLKINVX1 U954 ( .A(PC_4[30]), .Y(n561) );
  OAI22XL U955 ( .A0(n1380), .A1(n444), .B0(n439), .B1(n562), .Y(PC_4_w[29])
         );
  CLKINVX1 U956 ( .A(PC_4[29]), .Y(n562) );
  OAI22XL U957 ( .A0(n1381), .A1(n444), .B0(n439), .B1(n566), .Y(PC_4_w[28])
         );
  CLKINVX1 U958 ( .A(PC_4[28]), .Y(n566) );
  OAI22XL U959 ( .A0(n909), .A1(n451), .B0(n707), .B1(n437), .Y(inst_w[26]) );
  CLKINVX1 U960 ( .A(ICACHE_rdata[26]), .Y(n707) );
  OAI22XL U961 ( .A0(n1378), .A1(n444), .B0(n439), .B1(n556), .Y(PC_4_w[31])
         );
  CLKINVX1 U962 ( .A(PC_4[31]), .Y(n556) );
  OAI22XL U963 ( .A0(n1382), .A1(n448), .B0(n437), .B1(n644), .Y(PC_4_w[1]) );
  OAI22XL U964 ( .A0(n1383), .A1(n446), .B0(n441), .B1(n1579), .Y(PC_4_w[0])
         );
  OAI222XL U965 ( .A0(n1515), .A1(n255), .B0(n831), .B1(n256), .C0(n864), .C1(
        n250), .Y(n1377) );
  CLKINVX1 U966 ( .A(readreg1_forward[9]), .Y(n1515) );
  OAI222XL U967 ( .A0(n1519), .A1(n252), .B0(n829), .B1(n261), .C0(n862), .C1(
        n250), .Y(n1375) );
  CLKINVX1 U968 ( .A(readreg1_forward[7]), .Y(n1519) );
  NAND2X1 U969 ( .A(n548), .B(n549), .Y(PC_w[31]) );
  AOI222XL U970 ( .A0(N329), .A1(n242), .B0(PC_4[31]), .B1(n550), .C0(n245), 
        .C1(n551), .Y(n549) );
  AOI222XL U971 ( .A0(n236), .A1(ICACHE_addr[29]), .B0(N117), .B1(n233), .C0(
        n231), .C1(PC_4_r[31]), .Y(n548) );
  NAND2X1 U972 ( .A(n553), .B(n554), .Y(PC_w[30]) );
  AOI222XL U973 ( .A0(N328), .A1(n242), .B0(PC_4[30]), .B1(n550), .C0(n245), 
        .C1(n555), .Y(n554) );
  AOI222XL U974 ( .A0(n236), .A1(ICACHE_addr[28]), .B0(N116), .B1(n233), .C0(
        n231), .C1(PC_4_r[30]), .Y(n553) );
  NAND2X1 U975 ( .A(n563), .B(n564), .Y(PC_w[29]) );
  AOI222XL U976 ( .A0(N327), .A1(n242), .B0(PC_4[29]), .B1(n550), .C0(n245), 
        .C1(n565), .Y(n564) );
  AOI222XL U977 ( .A0(n236), .A1(ICACHE_addr[27]), .B0(N115), .B1(n233), .C0(
        n231), .C1(PC_4_r[29]), .Y(n563) );
  NAND2X1 U978 ( .A(n567), .B(n568), .Y(PC_w[28]) );
  AOI222XL U979 ( .A0(N326), .A1(n242), .B0(PC_4[28]), .B1(n550), .C0(n245), 
        .C1(n569), .Y(n568) );
  AOI222XL U980 ( .A0(n236), .A1(ICACHE_addr[26]), .B0(N114), .B1(n233), .C0(
        n231), .C1(PC_4_r[28]), .Y(n567) );
  NAND2X1 U981 ( .A(n622), .B(n623), .Y(PC_w[1]) );
  AOI222XL U982 ( .A0(n235), .A1(PC_r[1]), .B0(N87), .B1(n509), .C0(n232), 
        .C1(PC_4_r[1]), .Y(n622) );
  AOI222XL U983 ( .A0(N299), .A1(n242), .B0(PC_4[1]), .B1(n42), .C0(n245), 
        .C1(n625), .Y(n623) );
  NAND2X1 U984 ( .A(n690), .B(n691), .Y(PC_w[0]) );
  AOI222XL U985 ( .A0(n235), .A1(PC_r[0]), .B0(N86), .B1(n234), .C0(n231), 
        .C1(PC_4_r[0]), .Y(n690) );
  AOI222XL U986 ( .A0(N298), .A1(n242), .B0(PC_4[0]), .B1(n42), .C0(n245), 
        .C1(n692), .Y(n691) );
  NAND2X1 U987 ( .A(n645), .B(n646), .Y(PC_w[16]) );
  AOI222XL U988 ( .A0(n235), .A1(ICACHE_addr[14]), .B0(N102), .B1(n234), .C0(
        n232), .C1(PC_4_r[16]), .Y(n645) );
  AOI221XL U989 ( .A0(n244), .A1(n647), .B0(N314), .B1(n242), .C0(n648), .Y(
        n646) );
  NAND2X1 U990 ( .A(n651), .B(n652), .Y(PC_w[15]) );
  AOI222XL U991 ( .A0(n236), .A1(ICACHE_addr[13]), .B0(N101), .B1(n234), .C0(
        n231), .C1(PC_4_r[15]), .Y(n651) );
  AOI221XL U992 ( .A0(n245), .A1(n653), .B0(N313), .B1(n242), .C0(n654), .Y(
        n652) );
  NAND2X1 U993 ( .A(n663), .B(n664), .Y(PC_w[13]) );
  AOI222XL U994 ( .A0(n235), .A1(ICACHE_addr[11]), .B0(N99), .B1(n234), .C0(
        n232), .C1(PC_4_r[13]), .Y(n663) );
  AOI221XL U995 ( .A0(n244), .A1(n665), .B0(N311), .B1(n242), .C0(n666), .Y(
        n664) );
  NAND2X1 U996 ( .A(n669), .B(n670), .Y(PC_w[12]) );
  AOI222XL U997 ( .A0(n235), .A1(ICACHE_addr[10]), .B0(N98), .B1(n234), .C0(
        n231), .C1(PC_4_r[12]), .Y(n669) );
  AOI221XL U998 ( .A0(n245), .A1(n671), .B0(N310), .B1(n242), .C0(n672), .Y(
        n670) );
  NAND2X1 U999 ( .A(n675), .B(n676), .Y(PC_w[11]) );
  AOI222XL U1000 ( .A0(n235), .A1(ICACHE_addr[9]), .B0(N97), .B1(n234), .C0(
        n232), .C1(PC_4_r[11]), .Y(n675) );
  AOI221XL U1001 ( .A0(n501), .A1(n677), .B0(N309), .B1(n242), .C0(n678), .Y(
        n676) );
  NAND2X1 U1002 ( .A(n681), .B(n682), .Y(PC_w[10]) );
  AOI222XL U1003 ( .A0(n235), .A1(ICACHE_addr[8]), .B0(N96), .B1(n234), .C0(
        n231), .C1(PC_4_r[10]), .Y(n681) );
  AOI221XL U1004 ( .A0(n501), .A1(n683), .B0(N308), .B1(n242), .C0(n684), .Y(
        n682) );
  NAND2X1 U1005 ( .A(n499), .B(n500), .Y(PC_w[9]) );
  AOI222XL U1006 ( .A0(n235), .A1(ICACHE_addr[7]), .B0(N95), .B1(n233), .C0(
        n231), .C1(PC_4_r[9]), .Y(n499) );
  AOI221XL U1007 ( .A0(n244), .A1(n502), .B0(N307), .B1(n242), .C0(n504), .Y(
        n500) );
  NAND2X1 U1008 ( .A(n512), .B(n513), .Y(PC_w[8]) );
  AOI222XL U1009 ( .A0(n236), .A1(ICACHE_addr[6]), .B0(N94), .B1(n233), .C0(
        n231), .C1(PC_4_r[8]), .Y(n512) );
  AOI221XL U1010 ( .A0(n245), .A1(n514), .B0(N306), .B1(n243), .C0(n515), .Y(
        n513) );
  NAND2X1 U1011 ( .A(n518), .B(n519), .Y(PC_w[7]) );
  AOI222XL U1012 ( .A0(n236), .A1(ICACHE_addr[5]), .B0(N93), .B1(n233), .C0(
        n231), .C1(PC_4_r[7]), .Y(n518) );
  AOI221XL U1013 ( .A0(n245), .A1(n520), .B0(N305), .B1(n242), .C0(n521), .Y(
        n519) );
  NAND2X1 U1014 ( .A(n524), .B(n525), .Y(PC_w[6]) );
  AOI222XL U1015 ( .A0(n236), .A1(ICACHE_addr[4]), .B0(N92), .B1(n233), .C0(
        n231), .C1(PC_4_r[6]), .Y(n524) );
  AOI221XL U1016 ( .A0(n245), .A1(n526), .B0(N304), .B1(n243), .C0(n527), .Y(
        n525) );
  NAND2X1 U1017 ( .A(n530), .B(n531), .Y(PC_w[5]) );
  AOI222XL U1018 ( .A0(n236), .A1(ICACHE_addr[3]), .B0(N91), .B1(n233), .C0(
        n231), .C1(PC_4_r[5]), .Y(n530) );
  AOI221XL U1019 ( .A0(n245), .A1(n532), .B0(N303), .B1(n242), .C0(n533), .Y(
        n531) );
  NAND2X1 U1020 ( .A(n536), .B(n537), .Y(PC_w[4]) );
  AOI222XL U1021 ( .A0(n236), .A1(ICACHE_addr[2]), .B0(N90), .B1(n233), .C0(
        n231), .C1(PC_4_r[4]), .Y(n536) );
  AOI221XL U1022 ( .A0(n245), .A1(n538), .B0(N302), .B1(n243), .C0(n539), .Y(
        n537) );
  NAND2X1 U1023 ( .A(n542), .B(n543), .Y(PC_w[3]) );
  AOI222XL U1024 ( .A0(n236), .A1(ICACHE_addr[1]), .B0(N89), .B1(n233), .C0(
        n231), .C1(PC_4_r[3]), .Y(n542) );
  AOI221XL U1025 ( .A0(n245), .A1(n544), .B0(N301), .B1(n242), .C0(n545), .Y(
        n543) );
  OAI222XL U1026 ( .A0(n1505), .A1(n255), .B0(n805), .B1(n256), .C0(n838), 
        .C1(n250), .Y(n1351) );
  CLKINVX1 U1027 ( .A(readreg1_forward[14]), .Y(n1505) );
  OAI222XL U1028 ( .A0(n1517), .A1(n252), .B0(n830), .B1(n261), .C0(n863), 
        .C1(n250), .Y(n1376) );
  CLKINVX1 U1029 ( .A(readreg1_forward[8]), .Y(n1517) );
  OAI222XL U1030 ( .A0(n1509), .A1(n255), .B0(n803), .B1(n256), .C0(n836), 
        .C1(n250), .Y(n1349) );
  CLKINVX1 U1031 ( .A(readreg1_forward[12]), .Y(n1509) );
  OAI222XL U1032 ( .A0(n1511), .A1(n255), .B0(n802), .B1(n256), .C0(n835), 
        .C1(n251), .Y(n1348) );
  CLKINVX1 U1033 ( .A(readreg1_forward[11]), .Y(n1511) );
  OAI222XL U1034 ( .A0(n1507), .A1(n255), .B0(n804), .B1(n256), .C0(n837), 
        .C1(n251), .Y(n1350) );
  CLKINVX1 U1035 ( .A(readreg1_forward[13]), .Y(n1507) );
  OAI222XL U1036 ( .A0(n1513), .A1(n252), .B0(n801), .B1(n256), .C0(n834), 
        .C1(n251), .Y(n1347) );
  CLKINVX1 U1037 ( .A(readreg1_forward[10]), .Y(n1513) );
  CLKBUFX3 U1038 ( .A(n189), .Y(n295) );
  NOR2X1 U1039 ( .A(ICACHE_stall), .B(DCACHE_stall), .Y(n189) );
  OAI222XL U1040 ( .A0(n311), .A1(n1414), .B0(n293), .B1(n1048), .C0(n505), 
        .C1(n289), .Y(n1201) );
  CLKINVX1 U1041 ( .A(ALUresult[15]), .Y(n505) );
  OAI222XL U1042 ( .A0(n311), .A1(n1408), .B0(n293), .B1(n1036), .C0(n491), 
        .C1(n287), .Y(n1189) );
  CLKINVX1 U1043 ( .A(ALUresult[21]), .Y(n491) );
  OAI222XL U1044 ( .A0(n311), .A1(n1411), .B0(n293), .B1(n1042), .C0(n494), 
        .C1(n289), .Y(n1195) );
  CLKINVX1 U1045 ( .A(ALUresult[18]), .Y(n494) );
  OAI222XL U1046 ( .A0(n1485), .A1(n255), .B0(n816), .B1(n261), .C0(n849), 
        .C1(n250), .Y(n1362) );
  CLKINVX1 U1047 ( .A(readreg1_forward[24]), .Y(n1485) );
  OAI222XL U1048 ( .A0(n1411), .A1(n230), .B0(n415), .B1(n228), .C0(n1317), 
        .C1(n226), .Y(n726) );
  OAI222XL U1049 ( .A0(n1412), .A1(n230), .B0(n413), .B1(n228), .C0(n1319), 
        .C1(n226), .Y(n727) );
  OAI222XL U1050 ( .A0(n1413), .A1(n230), .B0(n411), .B1(n228), .C0(n1321), 
        .C1(n226), .Y(n728) );
  OAI222XL U1051 ( .A0(n1427), .A1(n229), .B0(n443), .B1(n228), .C0(n1465), 
        .C1(n225), .Y(n762) );
  OAI222XL U1052 ( .A0(n1428), .A1(n229), .B0(n420), .B1(n227), .C0(n1467), 
        .C1(n225), .Y(n763) );
  OAI222XL U1053 ( .A0(n1469), .A1(n226), .B0(n1429), .B1(n230), .C0(n396), 
        .C1(n227), .Y(n764) );
  OAI222XL U1054 ( .A0(n309), .A1(n1415), .B0(n293), .B1(n1050), .C0(n506), 
        .C1(n289), .Y(n1203) );
  CLKINVX1 U1055 ( .A(ALUresult[14]), .Y(n506) );
  OAI222XL U1056 ( .A0(n311), .A1(n1416), .B0(n293), .B1(n1052), .C0(n511), 
        .C1(n289), .Y(n1205) );
  CLKINVX1 U1057 ( .A(ALUresult[13]), .Y(n511) );
  OAI222XL U1058 ( .A0(n311), .A1(n1418), .B0(n293), .B1(n1056), .C0(n517), 
        .C1(n289), .Y(n1209) );
  CLKINVX1 U1059 ( .A(ALUresult[11]), .Y(n517) );
  OAI222XL U1060 ( .A0(n311), .A1(n1419), .B0(n291), .B1(n1058), .C0(n522), 
        .C1(n289), .Y(n1211) );
  CLKINVX1 U1061 ( .A(ALUresult[10]), .Y(n522) );
  OAI222XL U1062 ( .A0(n309), .A1(n1421), .B0(n291), .B1(n1062), .C0(n528), 
        .C1(n289), .Y(n1215) );
  CLKINVX1 U1063 ( .A(ALUresult[8]), .Y(n528) );
  OAI222XL U1064 ( .A0(n309), .A1(n1423), .B0(n291), .B1(n1066), .C0(n534), 
        .C1(n289), .Y(n1219) );
  CLKINVX1 U1065 ( .A(ALUresult[6]), .Y(n534) );
  OAI222XL U1066 ( .A0(n309), .A1(n1424), .B0(n291), .B1(n1068), .C0(n535), 
        .C1(n287), .Y(n1221) );
  CLKINVX1 U1067 ( .A(ALUresult[5]), .Y(n535) );
  OAI222XL U1068 ( .A0(n309), .A1(n1426), .B0(n291), .B1(n1072), .C0(n541), 
        .C1(n289), .Y(n1225) );
  CLKINVX1 U1069 ( .A(ALUresult[3]), .Y(n541) );
  OAI222XL U1070 ( .A0(n309), .A1(n1427), .B0(n291), .B1(n1074), .C0(n546), 
        .C1(n223), .Y(n1227) );
  CLKINVX1 U1071 ( .A(ALUresult[2]), .Y(n546) );
  OAI222XL U1072 ( .A0(n1393), .A1(n253), .B0(n1078), .B1(n254), .C0(n1079), 
        .C1(n309), .Y(n1231) );
  OAI222XL U1073 ( .A0(n1392), .A1(n253), .B0(n1081), .B1(n254), .C0(n1082), 
        .C1(n309), .Y(n1233) );
  OAI222XL U1074 ( .A0(n1391), .A1(n253), .B0(n1084), .B1(n254), .C0(n1085), 
        .C1(n309), .Y(n1235) );
  OAI222XL U1075 ( .A0(n1390), .A1(n253), .B0(n1395), .B1(n254), .C0(n1087), 
        .C1(n307), .Y(n1237) );
  OAI222XL U1076 ( .A0(n1394), .A1(n253), .B0(n1089), .B1(n254), .C0(n1091), 
        .C1(n307), .Y(n1239) );
  OAI221XL U1077 ( .A0(n1388), .A1(n408), .B0(n1394), .B1(n387), .C0(n498), 
        .Y(RegRt_idex_w[0]) );
  OAI221XL U1078 ( .A0(n1387), .A1(n402), .B0(n1393), .B1(n385), .C0(n498), 
        .Y(RegRt_idex_w[1]) );
  OAI221XL U1079 ( .A0(n1386), .A1(n404), .B0(n1392), .B1(n385), .C0(n498), 
        .Y(RegRt_idex_w[2]) );
  OAI221XL U1080 ( .A0(n1385), .A1(n400), .B0(n1391), .B1(n387), .C0(n498), 
        .Y(RegRt_idex_w[3]) );
  OAI221XL U1081 ( .A0(n1384), .A1(n433), .B0(n1390), .B1(n387), .C0(n498), 
        .Y(RegRt_idex_w[4]) );
  XOR2X1 U1082 ( .A(n629), .B(n719), .Y(n718) );
  OAI222XL U1083 ( .A0(n1410), .A1(n229), .B0(n417), .B1(n227), .C0(n1315), 
        .C1(n225), .Y(n719) );
  XOR2X1 U1084 ( .A(n551), .B(n749), .Y(n748) );
  OAI222XL U1085 ( .A0(n1398), .A1(n230), .B0(n447), .B1(n228), .C0(n1291), 
        .C1(n225), .Y(n749) );
  XOR2X1 U1086 ( .A(n600), .B(n733), .Y(n732) );
  OAI222XL U1087 ( .A0(n1406), .A1(n230), .B0(n428), .B1(n228), .C0(n1307), 
        .C1(n226), .Y(n733) );
  XOR2X1 U1088 ( .A(n576), .B(n741), .Y(n740) );
  OAI222XL U1089 ( .A0(n1402), .A1(n230), .B0(n436), .B1(n228), .C0(n1299), 
        .C1(n226), .Y(n741) );
  XOR2X1 U1090 ( .A(n544), .B(n761), .Y(n760) );
  OAI222XL U1091 ( .A0(n1426), .A1(n230), .B0(n450), .B1(n228), .C0(n1463), 
        .C1(n225), .Y(n761) );
  XOR2X1 U1092 ( .A(n520), .B(n769), .Y(n768) );
  OAI222XL U1093 ( .A0(n1422), .A1(n229), .B0(n459), .B1(n227), .C0(n1339), 
        .C1(n226), .Y(n769) );
  XOR2X1 U1094 ( .A(n677), .B(n777), .Y(n776) );
  OAI222XL U1095 ( .A0(n1418), .A1(n230), .B0(n401), .B1(n228), .C0(n1331), 
        .C1(n226), .Y(n777) );
  XOR2X1 U1096 ( .A(n653), .B(n785), .Y(n784) );
  OAI222XL U1097 ( .A0(n1414), .A1(n229), .B0(n409), .B1(n227), .C0(n1323), 
        .C1(n226), .Y(n785) );
  XOR2X1 U1098 ( .A(n555), .B(n750), .Y(n747) );
  OAI222XL U1099 ( .A0(n1399), .A1(n230), .B0(n445), .B1(n228), .C0(n1293), 
        .C1(n225), .Y(n750) );
  XOR2X1 U1100 ( .A(n606), .B(n734), .Y(n731) );
  OAI222XL U1101 ( .A0(n1407), .A1(n230), .B0(n426), .B1(n228), .C0(n1309), 
        .C1(n226), .Y(n734) );
  XOR2X1 U1102 ( .A(n582), .B(n742), .Y(n739) );
  OAI222XL U1103 ( .A0(n1403), .A1(n230), .B0(n434), .B1(n228), .C0(n1301), 
        .C1(n225), .Y(n742) );
  XOR2X1 U1104 ( .A(n526), .B(n770), .Y(n767) );
  OAI222XL U1105 ( .A0(n1423), .A1(n229), .B0(n457), .B1(n227), .C0(n1341), 
        .C1(n226), .Y(n770) );
  XOR2X1 U1106 ( .A(n683), .B(n778), .Y(n775) );
  OAI222XL U1107 ( .A0(n1419), .A1(n229), .B0(n399), .B1(n227), .C0(n1333), 
        .C1(n225), .Y(n778) );
  XOR2X1 U1108 ( .A(n659), .B(n786), .Y(n783) );
  OAI222XL U1109 ( .A0(n1415), .A1(n229), .B0(n407), .B1(n227), .C0(n1325), 
        .C1(n226), .Y(n786) );
  XOR2X1 U1110 ( .A(n569), .B(n752), .Y(n745) );
  OAI222XL U1111 ( .A0(n1401), .A1(n230), .B0(n438), .B1(n228), .C0(n1297), 
        .C1(n225), .Y(n752) );
  XOR2X1 U1112 ( .A(n618), .B(n736), .Y(n729) );
  OAI222XL U1113 ( .A0(n1409), .A1(n230), .B0(n422), .B1(n228), .C0(n1313), 
        .C1(n225), .Y(n736) );
  XOR2X1 U1114 ( .A(n594), .B(n744), .Y(n737) );
  OAI222XL U1115 ( .A0(n1405), .A1(n230), .B0(n430), .B1(n228), .C0(n1305), 
        .C1(n225), .Y(n744) );
  XOR2X1 U1116 ( .A(n538), .B(n772), .Y(n765) );
  OAI222XL U1117 ( .A0(n1425), .A1(n229), .B0(n453), .B1(n227), .C0(n1345), 
        .C1(n722), .Y(n772) );
  XOR2X1 U1118 ( .A(n514), .B(n780), .Y(n773) );
  OAI222XL U1119 ( .A0(n1421), .A1(n229), .B0(n461), .B1(n227), .C0(n1337), 
        .C1(n722), .Y(n780) );
  XOR2X1 U1120 ( .A(n671), .B(n788), .Y(n781) );
  OAI222XL U1121 ( .A0(n1417), .A1(n229), .B0(n403), .B1(n227), .C0(n1329), 
        .C1(n225), .Y(n788) );
  XOR2X1 U1122 ( .A(n565), .B(n751), .Y(n746) );
  OAI222XL U1123 ( .A0(n1400), .A1(n230), .B0(n440), .B1(n228), .C0(n1295), 
        .C1(n225), .Y(n751) );
  XOR2X1 U1124 ( .A(n612), .B(n735), .Y(n730) );
  OAI222XL U1125 ( .A0(n1408), .A1(n230), .B0(n424), .B1(n228), .C0(n1311), 
        .C1(n226), .Y(n735) );
  XOR2X1 U1126 ( .A(n588), .B(n743), .Y(n738) );
  OAI222XL U1127 ( .A0(n1404), .A1(n230), .B0(n432), .B1(n228), .C0(n1303), 
        .C1(n225), .Y(n743) );
  XOR2X1 U1128 ( .A(n532), .B(n771), .Y(n766) );
  OAI222XL U1129 ( .A0(n1424), .A1(n229), .B0(n455), .B1(n227), .C0(n1343), 
        .C1(n722), .Y(n771) );
  XOR2X1 U1130 ( .A(n502), .B(n779), .Y(n774) );
  OAI222XL U1131 ( .A0(n1420), .A1(n229), .B0(n463), .B1(n227), .C0(n1335), 
        .C1(n722), .Y(n779) );
  XOR2X1 U1132 ( .A(n665), .B(n787), .Y(n782) );
  OAI222XL U1133 ( .A0(n1416), .A1(n229), .B0(n405), .B1(n227), .C0(n1327), 
        .C1(n226), .Y(n787) );
  NAND2X1 U1134 ( .A(n1090), .B(n387), .Y(n253) );
  OAI211X1 U1135 ( .A0(n696), .A1(n702), .B0(n1288), .C0(n1289), .Y(n695) );
  CLKINVX1 U1136 ( .A(n686), .Y(n702) );
  AOI32X1 U1137 ( .A0(take), .A1(n706), .A2(ICACHE_rdata[28]), .B0(
        ICACHE_rdata[27]), .B1(n705), .Y(n696) );
  NAND2X1 U1138 ( .A(taken), .B(take_r), .Y(n693) );
  OAI22XL U1139 ( .A0(n1078), .A1(n377), .B0(n398), .B1(n1574), .Y(
        RegRd_idex_w[1]) );
  OAI22XL U1140 ( .A0(n1081), .A1(n379), .B0(n398), .B1(n1572), .Y(
        RegRd_idex_w[2]) );
  OAI22XL U1141 ( .A0(n1084), .A1(n375), .B0(n398), .B1(n1570), .Y(
        RegRd_idex_w[3]) );
  OAI22XL U1142 ( .A0(n1089), .A1(n377), .B0(n398), .B1(n1536), .Y(
        RegRd_idex_w[0]) );
  OAI22XL U1143 ( .A0(n793), .A1(n387), .B0(n947), .B1(n412), .Y(
        Funct_idex_w[0]) );
  OAI22XL U1144 ( .A0(n379), .A1(n1578), .B0(n947), .B1(n406), .Y(
        sign_ext_w[0]) );
  OAI22XL U1145 ( .A0(n794), .A1(n387), .B0(n948), .B1(n414), .Y(
        Funct_idex_w[1]) );
  OAI22XL U1146 ( .A0(n379), .A1(n1552), .B0(n948), .B1(n402), .Y(
        sign_ext_w[1]) );
  OAI22XL U1147 ( .A0(n795), .A1(n387), .B0(n949), .B1(n414), .Y(
        Funct_idex_w[2]) );
  OAI22XL U1148 ( .A0(n379), .A1(n1551), .B0(n949), .B1(n423), .Y(
        sign_ext_w[2]) );
  OAI22XL U1149 ( .A0(n796), .A1(n387), .B0(n950), .B1(n412), .Y(
        Funct_idex_w[3]) );
  OAI22XL U1150 ( .A0(n379), .A1(n1549), .B0(n950), .B1(n423), .Y(
        sign_ext_w[3]) );
  OAI22XL U1151 ( .A0(n797), .A1(n387), .B0(n951), .B1(n412), .Y(
        Funct_idex_w[4]) );
  OAI22XL U1152 ( .A0(n379), .A1(n1548), .B0(n951), .B1(n423), .Y(
        sign_ext_w[4]) );
  OAI22XL U1153 ( .A0(n798), .A1(n387), .B0(n952), .B1(n412), .Y(
        Funct_idex_w[5]) );
  OAI22XL U1154 ( .A0(n379), .A1(n1547), .B0(n952), .B1(n423), .Y(
        sign_ext_w[5]) );
  OAI22XL U1155 ( .A0(n1103), .A1(n387), .B0(n1378), .B1(n421), .Y(
        PC_4_idex_w[31]) );
  OAI22XL U1156 ( .A0(n1018), .A1(n387), .B0(n1379), .B1(n421), .Y(
        PC_4_idex_w[30]) );
  OAI22XL U1157 ( .A0(n1020), .A1(n381), .B0(n1380), .B1(n418), .Y(
        PC_4_idex_w[29]) );
  OAI22XL U1158 ( .A0(n1022), .A1(n379), .B0(n1381), .B1(n418), .Y(
        PC_4_idex_w[28]) );
  OAI22XL U1159 ( .A0(n1024), .A1(n375), .B0(n889), .B1(n418), .Y(
        PC_4_idex_w[27]) );
  OAI22XL U1160 ( .A0(n1026), .A1(n383), .B0(n888), .B1(n418), .Y(
        PC_4_idex_w[26]) );
  OAI22XL U1161 ( .A0(n1028), .A1(n385), .B0(n887), .B1(n418), .Y(
        PC_4_idex_w[25]) );
  OAI22XL U1162 ( .A0(n1030), .A1(n385), .B0(n886), .B1(n418), .Y(
        PC_4_idex_w[24]) );
  OAI22XL U1163 ( .A0(n1032), .A1(n379), .B0(n885), .B1(n418), .Y(
        PC_4_idex_w[23]) );
  OAI22XL U1164 ( .A0(n1034), .A1(n373), .B0(n884), .B1(n418), .Y(
        PC_4_idex_w[22]) );
  OAI22XL U1165 ( .A0(n1036), .A1(n387), .B0(n883), .B1(n416), .Y(
        PC_4_idex_w[21]) );
  OAI22XL U1166 ( .A0(n1038), .A1(n385), .B0(n882), .B1(n416), .Y(
        PC_4_idex_w[20]) );
  OAI22XL U1167 ( .A0(n1040), .A1(n377), .B0(n881), .B1(n416), .Y(
        PC_4_idex_w[19]) );
  OAI22XL U1168 ( .A0(n1042), .A1(n375), .B0(n880), .B1(n418), .Y(
        PC_4_idex_w[18]) );
  OAI22XL U1169 ( .A0(n1044), .A1(n387), .B0(n879), .B1(n416), .Y(
        PC_4_idex_w[17]) );
  OAI22XL U1170 ( .A0(n1046), .A1(n385), .B0(n878), .B1(n416), .Y(
        PC_4_idex_w[16]) );
  OAI22XL U1171 ( .A0(n1048), .A1(n385), .B0(n877), .B1(n416), .Y(
        PC_4_idex_w[15]) );
  OAI22XL U1172 ( .A0(n1050), .A1(n385), .B0(n876), .B1(n416), .Y(
        PC_4_idex_w[14]) );
  OAI22XL U1173 ( .A0(n1052), .A1(n385), .B0(n875), .B1(n416), .Y(
        PC_4_idex_w[13]) );
  OAI22XL U1174 ( .A0(n1054), .A1(n385), .B0(n874), .B1(n414), .Y(
        PC_4_idex_w[12]) );
  OAI22XL U1175 ( .A0(n1056), .A1(n385), .B0(n873), .B1(n414), .Y(
        PC_4_idex_w[11]) );
  OAI22XL U1176 ( .A0(n1058), .A1(n385), .B0(n872), .B1(n414), .Y(
        PC_4_idex_w[10]) );
  OAI22XL U1177 ( .A0(n1060), .A1(n387), .B0(n897), .B1(n421), .Y(
        PC_4_idex_w[9]) );
  OAI22XL U1178 ( .A0(n1062), .A1(n381), .B0(n896), .B1(n421), .Y(
        PC_4_idex_w[8]) );
  OAI22XL U1179 ( .A0(n1064), .A1(n387), .B0(n895), .B1(n421), .Y(
        PC_4_idex_w[7]) );
  OAI22XL U1180 ( .A0(n1066), .A1(n371), .B0(n894), .B1(n421), .Y(
        PC_4_idex_w[6]) );
  OAI22XL U1181 ( .A0(n1068), .A1(n371), .B0(n893), .B1(n421), .Y(
        PC_4_idex_w[5]) );
  OAI22XL U1182 ( .A0(n1070), .A1(n371), .B0(n892), .B1(n421), .Y(
        PC_4_idex_w[4]) );
  OAI22XL U1183 ( .A0(n1072), .A1(n371), .B0(n891), .B1(n421), .Y(
        PC_4_idex_w[3]) );
  OAI22XL U1184 ( .A0(n1074), .A1(n371), .B0(n890), .B1(n418), .Y(
        PC_4_idex_w[2]) );
  OAI22XL U1185 ( .A0(n1076), .A1(n383), .B0(n1382), .B1(n421), .Y(
        PC_4_idex_w[1]) );
  OAI22XL U1186 ( .A0(n1101), .A1(n385), .B0(n1383), .B1(n414), .Y(
        PC_4_idex_w[0]) );
  OAI22XL U1187 ( .A0(n1104), .A1(n319), .B0(n211), .B1(n297), .Y(n1249) );
  OAI22XL U1188 ( .A0(n1094), .A1(n297), .B0(n1093), .B1(n404), .Y(n1241) );
  OAI22XL U1189 ( .A0(n1096), .A1(n297), .B0(n1095), .B1(n423), .Y(n1242) );
  OAI22XL U1190 ( .A0(n1098), .A1(n297), .B0(n1097), .B1(n408), .Y(n1243) );
  OAI22XL U1191 ( .A0(n1104), .A1(n297), .B0(n1099), .B1(n400), .Y(n1244) );
  OAI22XL U1192 ( .A0(n898), .A1(n375), .B0(n904), .B1(n423), .Y(
        RegRs_idex_w[0]) );
  OAI22XL U1193 ( .A0(n899), .A1(n379), .B0(n905), .B1(n423), .Y(
        RegRs_idex_w[1]) );
  OAI22XL U1194 ( .A0(n900), .A1(n377), .B0(n906), .B1(n423), .Y(
        RegRs_idex_w[2]) );
  OAI22XL U1195 ( .A0(n901), .A1(n383), .B0(n907), .B1(n423), .Y(
        RegRs_idex_w[3]) );
  OAI22XL U1196 ( .A0(n902), .A1(n381), .B0(n908), .B1(n423), .Y(
        RegRs_idex_w[4]) );
  OAI22XL U1197 ( .A0(n866), .A1(n387), .B0(n909), .B1(n414), .Y(
        Opcode_idex_w[0]) );
  OAI22XL U1198 ( .A0(n867), .A1(n385), .B0(n910), .B1(n414), .Y(
        Opcode_idex_w[1]) );
  OAI22XL U1199 ( .A0(n868), .A1(n383), .B0(n911), .B1(n414), .Y(
        Opcode_idex_w[2]) );
  OAI22XL U1200 ( .A0(n869), .A1(n385), .B0(n912), .B1(n414), .Y(
        Opcode_idex_w[3]) );
  OAI22XL U1201 ( .A0(n870), .A1(n385), .B0(n913), .B1(n416), .Y(
        Opcode_idex_w[4]) );
  OAI22XL U1202 ( .A0(n871), .A1(n385), .B0(n914), .B1(n416), .Y(
        Opcode_idex_w[5]) );
  OAI22XL U1203 ( .A0(n1401), .A1(n333), .B0(n1021), .B1(n303), .Y(n1174) );
  OAI22XL U1204 ( .A0(n1402), .A1(n333), .B0(n1023), .B1(n303), .Y(n1176) );
  OAI22XL U1205 ( .A0(n1403), .A1(n333), .B0(n1025), .B1(n301), .Y(n1178) );
  OAI22XL U1206 ( .A0(n1404), .A1(n331), .B0(n1027), .B1(n301), .Y(n1180) );
  OAI22XL U1207 ( .A0(n1405), .A1(n331), .B0(n1029), .B1(n301), .Y(n1182) );
  OAI22XL U1208 ( .A0(n1406), .A1(n331), .B0(n1031), .B1(n301), .Y(n1184) );
  OAI22XL U1209 ( .A0(n1407), .A1(n331), .B0(n1033), .B1(n301), .Y(n1186) );
  OAI22XL U1210 ( .A0(n1408), .A1(n329), .B0(n1035), .B1(n301), .Y(n1188) );
  OAI22XL U1211 ( .A0(n1409), .A1(n329), .B0(n1037), .B1(n301), .Y(n1190) );
  OAI22XL U1212 ( .A0(n1410), .A1(n329), .B0(n1039), .B1(n301), .Y(n1192) );
  OAI22XL U1213 ( .A0(n1411), .A1(n329), .B0(n1041), .B1(n301), .Y(n1194) );
  OAI22XL U1214 ( .A0(n1412), .A1(n327), .B0(n1043), .B1(n301), .Y(n1196) );
  OAI22XL U1215 ( .A0(n1413), .A1(n327), .B0(n1045), .B1(n301), .Y(n1198) );
  OAI22XL U1216 ( .A0(n1414), .A1(n327), .B0(n1047), .B1(n301), .Y(n1200) );
  OAI22XL U1217 ( .A0(n1415), .A1(n327), .B0(n1049), .B1(n301), .Y(n1202) );
  OAI22XL U1218 ( .A0(n1416), .A1(n325), .B0(n1051), .B1(n299), .Y(n1204) );
  OAI22XL U1219 ( .A0(n1417), .A1(n325), .B0(n1053), .B1(n299), .Y(n1206) );
  OAI22XL U1220 ( .A0(n1418), .A1(n325), .B0(n1055), .B1(n299), .Y(n1208) );
  OAI22XL U1221 ( .A0(n1419), .A1(n325), .B0(n1057), .B1(n299), .Y(n1210) );
  OAI22XL U1222 ( .A0(n1420), .A1(n323), .B0(n1059), .B1(n299), .Y(n1212) );
  OAI22XL U1223 ( .A0(n1421), .A1(n323), .B0(n1061), .B1(n299), .Y(n1214) );
  OAI22XL U1224 ( .A0(n1422), .A1(n323), .B0(n1063), .B1(n299), .Y(n1216) );
  OAI22XL U1226 ( .A0(n1423), .A1(n323), .B0(n1065), .B1(n299), .Y(n1218) );
  OAI22XL U1227 ( .A0(n1424), .A1(n347), .B0(n1067), .B1(n299), .Y(n1220) );
  OAI22XL U1228 ( .A0(n1425), .A1(n351), .B0(n1069), .B1(n299), .Y(n1222) );
  OAI22XL U1229 ( .A0(n1426), .A1(n347), .B0(n1071), .B1(n299), .Y(n1224) );
  OAI22XL U1230 ( .A0(n1427), .A1(n351), .B0(n1073), .B1(n299), .Y(n1226) );
  OAI22XL U1232 ( .A0(n1428), .A1(n349), .B0(n1075), .B1(n299), .Y(n1228) );
  OAI22XL U1233 ( .A0(n1429), .A1(n321), .B0(n1100), .B1(n297), .Y(n1245) );
  OAI22XL U1234 ( .A0(n1532), .A1(n319), .B0(n954), .B1(n303), .Y(n1138) );
  OAI22XL U1235 ( .A0(n1502), .A1(n337), .B0(n988), .B1(n307), .Y(n1155) );
  OAI22XL U1236 ( .A0(n1398), .A1(n319), .B0(n1102), .B1(n297), .Y(n1247) );
  OAI22XL U1238 ( .A0(n1504), .A1(n333), .B0(n990), .B1(n307), .Y(n1156) );
  OAI22XL U1239 ( .A0(n1506), .A1(n337), .B0(n992), .B1(n307), .Y(n1157) );
  OAI22XL U1240 ( .A0(n1508), .A1(n337), .B0(n994), .B1(n307), .Y(n1158) );
  OAI22XL U1241 ( .A0(n1510), .A1(n337), .B0(n996), .B1(n307), .Y(n1159) );
  OAI22XL U1242 ( .A0(n1512), .A1(n335), .B0(n998), .B1(n307), .Y(n1160) );
  OAI22XL U1243 ( .A0(n1514), .A1(n335), .B0(n1000), .B1(n307), .Y(n1161) );
  OAI22XL U1244 ( .A0(n1516), .A1(n335), .B0(n1002), .B1(n305), .Y(n1162) );
  OAI22XL U1245 ( .A0(n1518), .A1(n335), .B0(n1004), .B1(n305), .Y(n1163) );
  OAI22XL U1246 ( .A0(n1520), .A1(n337), .B0(n1006), .B1(n305), .Y(n1164) );
  OAI22XL U1247 ( .A0(n1522), .A1(n335), .B0(n1008), .B1(n305), .Y(n1165) );
  OAI22XL U1248 ( .A0(n1524), .A1(n337), .B0(n1010), .B1(n305), .Y(n1166) );
  OAI22XL U1249 ( .A0(n1526), .A1(n335), .B0(n1012), .B1(n305), .Y(n1167) );
  OAI22XL U1250 ( .A0(n1528), .A1(n321), .B0(n1014), .B1(n305), .Y(n1168) );
  OAI22XL U1251 ( .A0(n1530), .A1(n349), .B0(n1016), .B1(n305), .Y(n1169) );
  OAI22XL U1252 ( .A0(n1399), .A1(n321), .B0(n1017), .B1(n303), .Y(n1170) );
  OAI22XL U1253 ( .A0(n1400), .A1(n349), .B0(n1019), .B1(n303), .Y(n1172) );
  OAI22XL U1254 ( .A0(n1079), .A1(n321), .B0(n1077), .B1(n297), .Y(n1230) );
  OAI22XL U1255 ( .A0(n1082), .A1(n321), .B0(n1080), .B1(n297), .Y(n1232) );
  OAI22XL U1256 ( .A0(n1085), .A1(n321), .B0(n1083), .B1(n297), .Y(n1234) );
  OAI22XL U1257 ( .A0(n1087), .A1(n321), .B0(n1086), .B1(n297), .Y(n1236) );
  OAI22XL U1258 ( .A0(n1091), .A1(n321), .B0(n1088), .B1(n297), .Y(n1238) );
  OAI22XL U1259 ( .A0(n1094), .A1(n321), .B0(n1092), .B1(n297), .Y(n1240) );
  OAI222XL U1260 ( .A0(n1499), .A1(n255), .B0(n808), .B1(n261), .C0(n841), 
        .C1(n250), .Y(n1354) );
  CLKINVX1 U1262 ( .A(readreg1_forward[17]), .Y(n1499) );
  OAI222XL U1263 ( .A0(n1497), .A1(n255), .B0(n809), .B1(n261), .C0(n842), 
        .C1(n250), .Y(n1355) );
  CLKINVX1 U1264 ( .A(readreg1_forward[18]), .Y(n1497) );
  OAI222XL U1265 ( .A0(n1487), .A1(n255), .B0(n815), .B1(n261), .C0(n848), 
        .C1(n251), .Y(n1361) );
  CLKINVX1 U1266 ( .A(readreg1_forward[23]), .Y(n1487) );
  OAI222XL U1267 ( .A0(n1503), .A1(n255), .B0(n806), .B1(n256), .C0(n839), 
        .C1(n250), .Y(n1352) );
  CLKINVX1 U1268 ( .A(readreg1_forward[15]), .Y(n1503) );
  OAI222XL U1269 ( .A0(n1501), .A1(n255), .B0(n807), .B1(n256), .C0(n840), 
        .C1(n250), .Y(n1353) );
  CLKINVX1 U1270 ( .A(readreg1_forward[16]), .Y(n1501) );
  OAI222XL U1271 ( .A0(n1471), .A1(n252), .B0(n824), .B1(n261), .C0(n857), 
        .C1(n250), .Y(n1370) );
  CLKINVX1 U1272 ( .A(readreg1_forward[31]), .Y(n1471) );
  OAI222XL U1273 ( .A0(n309), .A1(n1428), .B0(n291), .B1(n1076), .C0(n547), 
        .C1(n223), .Y(n1229) );
  CLKINVX1 U1274 ( .A(ALUresult[1]), .Y(n547) );
  OAI222XL U1275 ( .A0(n309), .A1(n1422), .B0(n291), .B1(n1064), .C0(n529), 
        .C1(n289), .Y(n1217) );
  CLKINVX1 U1276 ( .A(ALUresult[7]), .Y(n529) );
  OAI222XL U1277 ( .A0(n311), .A1(n1417), .B0(n293), .B1(n1054), .C0(n516), 
        .C1(n289), .Y(n1207) );
  CLKINVX1 U1278 ( .A(ALUresult[12]), .Y(n516) );
  OR2X1 U1279 ( .A(n1090), .B(n412), .Y(n254) );
  OAI2BB2XL U1280 ( .B0(n373), .B1(n903), .A0N(Shift), .A1N(n196), .Y(
        Shift_idex_w) );
  OAI2BB2XL U1281 ( .B0(n377), .B1(n799), .A0N(HI), .A1N(n196), .Y(HI_idex_w)
         );
  OAI2BB2XL U1282 ( .B0(n373), .B1(n832), .A0N(LO), .A1N(n196), .Y(LO_idex_w)
         );
  OAI2BB2XL U1283 ( .B0(n406), .B1(n1576), .A0N(n425), .A1N(shamt_idex_r[4]), 
        .Y(shamt_idex_w[4]) );
  OAI2BB2XL U1284 ( .B0(n392), .B1(n1545), .A0N(n425), .A1N(shamt_idex_r[0]), 
        .Y(shamt_idex_w[0]) );
  OAI2BB2XL U1286 ( .B0(n397), .B1(n1543), .A0N(n425), .A1N(shamt_idex_r[1]), 
        .Y(shamt_idex_w[1]) );
  OAI2BB2XL U1287 ( .B0(n397), .B1(n1541), .A0N(n425), .A1N(shamt_idex_r[2]), 
        .Y(shamt_idex_w[2]) );
  OAI2BB2XL U1288 ( .B0(n425), .B1(n1539), .A0N(n425), .A1N(shamt_idex_r[3]), 
        .Y(shamt_idex_w[3]) );
  OAI2BB2XL U1289 ( .B0(n373), .B1(n1090), .A0N(RegDst), .A1N(n196), .Y(
        RegDst_idex_w) );
  OAI2BB2XL U1290 ( .B0(n385), .B1(n1396), .A0N(Jump), .A1N(n196), .Y(
        Jump_idex_w) );
  OAI2BB2XL U1292 ( .B0(n373), .B1(n1397), .A0N(Div), .A1N(n196), .Y(
        Div_idex_w) );
  OAI2BB2XL U1293 ( .B0(n385), .B1(n865), .A0N(Mul), .A1N(n196), .Y(Mul_idex_w) );
  OAI2BB2XL U1294 ( .B0(n373), .B1(n1093), .A0N(RegWrite), .A1N(n196), .Y(
        RegWrite_idex_w) );
  OAI2BB2XL U1295 ( .B0(n379), .B1(n1095), .A0N(MemWrite), .A1N(n196), .Y(
        MemWrite_idex_w) );
  OAI2BB2XL U1296 ( .B0(n385), .B1(n1097), .A0N(MemRead), .A1N(n196), .Y(
        MemRead_idex_w) );
  OAI2BB2XL U1298 ( .B0(n373), .B1(n1099), .A0N(MemtoReg), .A1N(n196), .Y(
        MemtoReg_idex_w) );
  OAI21XL U1299 ( .A0(n1395), .A1(n381), .B0(n197), .Y(RegRd_idex_w[4]) );
  OAI222XL U1300 ( .A0(n309), .A1(n1429), .B0(n291), .B1(n1101), .C0(n552), 
        .C1(n223), .Y(n1246) );
  CLKINVX1 U1301 ( .A(ALUresult[0]), .Y(n552) );
  OAI222XL U1302 ( .A0(n1473), .A1(n252), .B0(n823), .B1(n261), .C0(n856), 
        .C1(n250), .Y(n1369) );
  CLKINVX1 U1303 ( .A(readreg1_forward[30]), .Y(n1473) );
  OAI222XL U1304 ( .A0(n1481), .A1(n255), .B0(n818), .B1(n261), .C0(n851), 
        .C1(n250), .Y(n1364) );
  CLKINVX1 U1305 ( .A(readreg1_forward[26]), .Y(n1481) );
  OAI222XL U1306 ( .A0(n1483), .A1(n255), .B0(n817), .B1(n261), .C0(n850), 
        .C1(n250), .Y(n1363) );
  CLKINVX1 U1307 ( .A(readreg1_forward[25]), .Y(n1483) );
  OAI222XL U1308 ( .A0(n1479), .A1(n255), .B0(n819), .B1(n261), .C0(n852), 
        .C1(n250), .Y(n1365) );
  CLKINVX1 U1310 ( .A(readreg1_forward[27]), .Y(n1479) );
  OAI222XL U1311 ( .A0(n1489), .A1(n255), .B0(n814), .B1(n261), .C0(n847), 
        .C1(n251), .Y(n1360) );
  CLKINVX1 U1312 ( .A(readreg1_forward[22]), .Y(n1489) );
  OAI222XL U1313 ( .A0(n1493), .A1(n255), .B0(n812), .B1(n261), .C0(n845), 
        .C1(n250), .Y(n1358) );
  CLKINVX1 U1314 ( .A(readreg1_forward[20]), .Y(n1493) );
  OAI222XL U1315 ( .A0(n1491), .A1(n255), .B0(n813), .B1(n261), .C0(n846), 
        .C1(n251), .Y(n1359) );
  CLKINVX1 U1316 ( .A(readreg1_forward[21]), .Y(n1491) );
  OAI222XL U1317 ( .A0(n1495), .A1(n255), .B0(n810), .B1(n261), .C0(n843), 
        .C1(n250), .Y(n1356) );
  CLKINVX1 U1318 ( .A(readreg1_forward[19]), .Y(n1495) );
  OAI222XL U1319 ( .A0(n1477), .A1(n255), .B0(n820), .B1(n261), .C0(n853), 
        .C1(n250), .Y(n1366) );
  CLKINVX1 U1320 ( .A(readreg1_forward[28]), .Y(n1477) );
  OAI222XL U1322 ( .A0(n1475), .A1(n252), .B0(n821), .B1(n261), .C0(n854), 
        .C1(n250), .Y(n1367) );
  CLKINVX1 U1323 ( .A(readreg1_forward[29]), .Y(n1475) );
  AO22X1 U1324 ( .A0(n400), .A1(ALUOp_idex_r[1]), .B0(ALUOp[1]), .B1(n196), 
        .Y(ALUOp_idex_w[1]) );
  AO22X1 U1325 ( .A0(n425), .A1(ALUOp_idex_r[0]), .B0(ALUOp[0]), .B1(n196), 
        .Y(ALUOp_idex_w[0]) );
  AO22X1 U1326 ( .A0(n321), .A1(n1106), .B0(DCACHE_rdata[0]), .B1(n313), .Y(
        n1250) );
  AO22X1 U1327 ( .A0(n351), .A1(n1107), .B0(DCACHE_rdata[1]), .B1(n313), .Y(
        n1251) );
  AO22X1 U1328 ( .A0(n351), .A1(n1108), .B0(DCACHE_rdata[2]), .B1(n313), .Y(
        n1252) );
  AO22X1 U1329 ( .A0(n347), .A1(n1109), .B0(DCACHE_rdata[3]), .B1(n313), .Y(
        n1253) );
  AO22X1 U1330 ( .A0(n321), .A1(n1110), .B0(DCACHE_rdata[4]), .B1(n313), .Y(
        n1254) );
  AO22X1 U1331 ( .A0(n317), .A1(n1111), .B0(DCACHE_rdata[5]), .B1(n313), .Y(
        n1255) );
  AO22X1 U1332 ( .A0(n349), .A1(n1112), .B0(DCACHE_rdata[6]), .B1(n315), .Y(
        n1256) );
  AO22X1 U1334 ( .A0(n347), .A1(n1113), .B0(DCACHE_rdata[7]), .B1(n313), .Y(
        n1257) );
  AO22X1 U1335 ( .A0(n351), .A1(n1114), .B0(DCACHE_rdata[8]), .B1(n313), .Y(
        n1258) );
  AO22X1 U1336 ( .A0(n321), .A1(n1115), .B0(DCACHE_rdata[9]), .B1(n313), .Y(
        n1259) );
  AO22X1 U1337 ( .A0(n351), .A1(n1116), .B0(DCACHE_rdata[10]), .B1(n313), .Y(
        n1260) );
  AO22X1 U1338 ( .A0(n345), .A1(n1117), .B0(DCACHE_rdata[11]), .B1(n313), .Y(
        n1261) );
  AO22X1 U1339 ( .A0(n345), .A1(n1118), .B0(DCACHE_rdata[12]), .B1(n313), .Y(
        n1262) );
  AO22X1 U1340 ( .A0(n345), .A1(n1119), .B0(DCACHE_rdata[13]), .B1(n313), .Y(
        n1263) );
  AO22X1 U1341 ( .A0(n345), .A1(n1120), .B0(DCACHE_rdata[14]), .B1(n313), .Y(
        n1264) );
  AO22X1 U1342 ( .A0(n345), .A1(n1121), .B0(DCACHE_rdata[15]), .B1(n313), .Y(
        n1265) );
  AO22X1 U1343 ( .A0(n347), .A1(n1122), .B0(DCACHE_rdata[16]), .B1(n315), .Y(
        n1266) );
  AO22X1 U1344 ( .A0(n347), .A1(n1123), .B0(DCACHE_rdata[17]), .B1(n315), .Y(
        n1267) );
  AO22X1 U1346 ( .A0(n347), .A1(n1124), .B0(DCACHE_rdata[18]), .B1(n315), .Y(
        n1268) );
  AO22X1 U1347 ( .A0(n347), .A1(n1125), .B0(DCACHE_rdata[19]), .B1(n315), .Y(
        n1269) );
  AO22X1 U1348 ( .A0(n347), .A1(n1126), .B0(DCACHE_rdata[20]), .B1(n315), .Y(
        n1270) );
  AO22X1 U1349 ( .A0(n347), .A1(n1127), .B0(DCACHE_rdata[21]), .B1(n315), .Y(
        n1271) );
  AO22X1 U1350 ( .A0(n349), .A1(n1128), .B0(DCACHE_rdata[22]), .B1(n315), .Y(
        n1272) );
  AO22X1 U1352 ( .A0(n349), .A1(n1129), .B0(DCACHE_rdata[23]), .B1(n315), .Y(
        n1273) );
  AO22X1 U1353 ( .A0(n349), .A1(n1130), .B0(DCACHE_rdata[24]), .B1(n315), .Y(
        n1274) );
  AO22X1 U1354 ( .A0(n349), .A1(n1131), .B0(DCACHE_rdata[25]), .B1(n315), .Y(
        n1275) );
  AO22X1 U1355 ( .A0(n349), .A1(n1132), .B0(DCACHE_rdata[26]), .B1(n315), .Y(
        n1276) );
  AO22X1 U1356 ( .A0(n349), .A1(n1133), .B0(DCACHE_rdata[27]), .B1(n315), .Y(
        n1277) );
  AO22X1 U1357 ( .A0(n351), .A1(n1134), .B0(DCACHE_rdata[28]), .B1(n315), .Y(
        n1278) );
  AO22X1 U1358 ( .A0(n351), .A1(n1135), .B0(DCACHE_rdata[29]), .B1(n315), .Y(
        n1279) );
  AO22X1 U1359 ( .A0(n351), .A1(n1136), .B0(DCACHE_rdata[30]), .B1(n315), .Y(
        n1280) );
  AO22X1 U1360 ( .A0(n351), .A1(n1137), .B0(DCACHE_rdata[31]), .B1(n313), .Y(
        n1281) );
  NOR2X1 U1361 ( .A(n709), .B(n710), .Y(N346) );
  OAI222XL U1362 ( .A0(n309), .A1(n1425), .B0(n291), .B1(n1070), .C0(n540), 
        .C1(n223), .Y(n1223) );
  CLKINVX1 U1363 ( .A(ALUresult[4]), .Y(n540) );
  OAI222XL U1364 ( .A0(n309), .A1(n1420), .B0(n291), .B1(n1060), .C0(n523), 
        .C1(n289), .Y(n1213) );
  CLKINVX1 U1365 ( .A(ALUresult[9]), .Y(n523) );
  CLKINVX1 U1366 ( .A(n372), .Y(n928) );
  AOI222XL U1367 ( .A0(LO_mul[31]), .A1(n279), .B0(LO_div[31]), .B1(n277), 
        .C0(n269), .C1(n46), .Y(n372) );
  OAI22XL U1368 ( .A0(n1472), .A1(n343), .B0(n956), .B1(n303), .Y(n1139) );
  OAI22XL U1369 ( .A0(n456), .A1(n343), .B0(n958), .B1(n303), .Y(n1140) );
  OAI22XL U1370 ( .A0(n1474), .A1(n343), .B0(n960), .B1(n303), .Y(n1141) );
  OAI22XL U1371 ( .A0(n1476), .A1(n343), .B0(n962), .B1(n303), .Y(n1142) );
  OAI22XL U1372 ( .A0(n1478), .A1(n341), .B0(n964), .B1(n303), .Y(n1143) );
  OAI22XL U1373 ( .A0(n1480), .A1(n341), .B0(n966), .B1(n303), .Y(n1144) );
  OAI22XL U1374 ( .A0(n1482), .A1(n341), .B0(n968), .B1(n303), .Y(n1145) );
  OAI22XL U1376 ( .A0(n1484), .A1(n341), .B0(n970), .B1(n305), .Y(n1146) );
  OAI22XL U1377 ( .A0(n1486), .A1(n339), .B0(n972), .B1(n305), .Y(n1147) );
  OAI22XL U1378 ( .A0(n1488), .A1(n339), .B0(n974), .B1(n305), .Y(n1148) );
  OAI22XL U1379 ( .A0(n1490), .A1(n339), .B0(n976), .B1(n305), .Y(n1149) );
  OAI22XL U1380 ( .A0(n1492), .A1(n339), .B0(n978), .B1(n305), .Y(n1150) );
  OAI22XL U1381 ( .A0(n1494), .A1(n341), .B0(n980), .B1(n307), .Y(n1151) );
  OAI22XL U1382 ( .A0(n1496), .A1(n339), .B0(n982), .B1(n307), .Y(n1152) );
  OAI22XL U1383 ( .A0(n1498), .A1(n343), .B0(n984), .B1(n307), .Y(n1153) );
  OAI22XL U1384 ( .A0(n1500), .A1(n343), .B0(n986), .B1(n303), .Y(n1154) );
  CLKINVX1 U1385 ( .A(n370), .Y(n929) );
  AOI222XL U1386 ( .A0(LO_mul[30]), .A1(n279), .B0(LO_div[30]), .B1(n277), 
        .C0(n269), .C1(n47), .Y(n370) );
  CLKINVX1 U1388 ( .A(n366), .Y(n931) );
  AOI222XL U1389 ( .A0(LO_mul[29]), .A1(n279), .B0(LO_div[29]), .B1(n277), 
        .C0(n269), .C1(n48), .Y(n366) );
  CLKINVX1 U1390 ( .A(n364), .Y(n932) );
  AOI222XL U1391 ( .A0(LO_mul[28]), .A1(n279), .B0(LO_div[28]), .B1(n277), 
        .C0(n269), .C1(n49), .Y(n364) );
  CLKINVX1 U1392 ( .A(n362), .Y(n933) );
  AOI222XL U1394 ( .A0(LO_mul[27]), .A1(n279), .B0(LO_div[27]), .B1(n277), 
        .C0(n269), .C1(n50), .Y(n362) );
  CLKINVX1 U1395 ( .A(n360), .Y(n934) );
  AOI222XL U1396 ( .A0(LO_mul[26]), .A1(n279), .B0(LO_div[26]), .B1(n277), 
        .C0(n269), .C1(n51), .Y(n360) );
  CLKINVX1 U1397 ( .A(n358), .Y(n935) );
  AOI222XL U1398 ( .A0(LO_mul[25]), .A1(n281), .B0(LO_div[25]), .B1(n277), 
        .C0(n269), .C1(n52), .Y(n358) );
  CLKINVX1 U1400 ( .A(n356), .Y(n936) );
  AOI222XL U1401 ( .A0(LO_mul[24]), .A1(n281), .B0(LO_div[24]), .B1(n277), 
        .C0(n269), .C1(n53), .Y(n356) );
  CLKINVX1 U1402 ( .A(n354), .Y(n937) );
  AOI222XL U1403 ( .A0(LO_mul[23]), .A1(n281), .B0(LO_div[23]), .B1(n275), 
        .C0(n267), .C1(n54), .Y(n354) );
  CLKINVX1 U1404 ( .A(n308), .Y(n979) );
  AOI222XL U1406 ( .A0(HI_mul[31]), .A1(n283), .B0(HI_div[31]), .B1(n271), 
        .C0(n263), .C1(n58), .Y(n308) );
  CLKINVX1 U1407 ( .A(n306), .Y(n981) );
  AOI222XL U1408 ( .A0(HI_mul[30]), .A1(n283), .B0(HI_div[30]), .B1(n273), 
        .C0(n267), .C1(n59), .Y(n306) );
  CLKINVX1 U1409 ( .A(n302), .Y(n985) );
  AOI222XL U1410 ( .A0(HI_mul[29]), .A1(n283), .B0(HI_div[29]), .B1(n273), 
        .C0(n265), .C1(n60), .Y(n302) );
  CLKINVX1 U1411 ( .A(n300), .Y(n987) );
  AOI222XL U1412 ( .A0(HI_mul[28]), .A1(n283), .B0(HI_div[28]), .B1(n273), 
        .C0(n267), .C1(n61), .Y(n300) );
  CLKINVX1 U1413 ( .A(n298), .Y(n989) );
  AOI222XL U1414 ( .A0(HI_mul[27]), .A1(n283), .B0(HI_div[27]), .B1(n273), 
        .C0(n263), .C1(n62), .Y(n298) );
  CLKINVX1 U1415 ( .A(n296), .Y(n991) );
  AOI222XL U1416 ( .A0(HI_mul[26]), .A1(n283), .B0(HI_div[26]), .B1(n273), 
        .C0(n265), .C1(n63), .Y(n296) );
  CLKINVX1 U1417 ( .A(n294), .Y(n993) );
  AOI222XL U1418 ( .A0(HI_mul[25]), .A1(n285), .B0(HI_div[25]), .B1(n273), 
        .C0(n260), .C1(n64), .Y(n294) );
  CLKINVX1 U1419 ( .A(n292), .Y(n995) );
  AOI222XL U1420 ( .A0(HI_mul[24]), .A1(n285), .B0(HI_div[24]), .B1(n273), 
        .C0(n260), .C1(n65), .Y(n292) );
  CLKINVX1 U1421 ( .A(n290), .Y(n997) );
  AOI222XL U1422 ( .A0(HI_mul[23]), .A1(n285), .B0(HI_div[23]), .B1(n273), 
        .C0(n260), .C1(n66), .Y(n290) );
  CLKINVX1 U1423 ( .A(n288), .Y(n999) );
  AOI222XL U1424 ( .A0(HI_mul[22]), .A1(n285), .B0(HI_div[22]), .B1(n273), 
        .C0(n260), .C1(n67), .Y(n288) );
  CLKINVX1 U1425 ( .A(n352), .Y(n938) );
  AOI222XL U1426 ( .A0(LO_mul[22]), .A1(n281), .B0(LO_div[22]), .B1(n275), 
        .C0(n267), .C1(n55), .Y(n352) );
  CLKINVX1 U1427 ( .A(n350), .Y(n939) );
  AOI222XL U1428 ( .A0(LO_mul[21]), .A1(n281), .B0(LO_div[21]), .B1(n275), 
        .C0(n267), .C1(n56), .Y(n350) );
  CLKINVX1 U1429 ( .A(n348), .Y(n940) );
  AOI222XL U1430 ( .A0(LO_mul[20]), .A1(n281), .B0(LO_div[20]), .B1(n275), 
        .C0(n267), .C1(n57), .Y(n348) );
  CLKINVX1 U1431 ( .A(n344), .Y(n942) );
  AOI222XL U1432 ( .A0(LO_mul[19]), .A1(n281), .B0(LO_div[19]), .B1(n275), 
        .C0(n267), .C1(n1663), .Y(n344) );
  CLKINVX1 U1433 ( .A(n342), .Y(n943) );
  AOI222XL U1434 ( .A0(LO_mul[18]), .A1(n281), .B0(LO_div[18]), .B1(n275), 
        .C0(n267), .C1(n1662), .Y(n342) );
  CLKINVX1 U1435 ( .A(n340), .Y(n944) );
  AOI222XL U1436 ( .A0(LO_mul[17]), .A1(n281), .B0(LO_div[17]), .B1(n275), 
        .C0(n267), .C1(n1661), .Y(n340) );
  CLKINVX1 U1437 ( .A(n338), .Y(n945) );
  AOI222XL U1438 ( .A0(LO_mul[16]), .A1(n281), .B0(LO_div[16]), .B1(n275), 
        .C0(n267), .C1(n1660), .Y(n338) );
  CLKINVX1 U1439 ( .A(n336), .Y(n946) );
  AOI222XL U1440 ( .A0(LO_mul[15]), .A1(n281), .B0(LO_div[15]), .B1(n275), 
        .C0(n267), .C1(n1659), .Y(n336) );
  CLKINVX1 U1441 ( .A(n334), .Y(n953) );
  AOI222XL U1442 ( .A0(LO_mul[14]), .A1(n281), .B0(LO_div[14]), .B1(n275), 
        .C0(n267), .C1(n1658), .Y(n334) );
  CLKINVX1 U1443 ( .A(n332), .Y(n955) );
  AOI222XL U1444 ( .A0(LO_mul[13]), .A1(n281), .B0(LO_div[13]), .B1(n275), 
        .C0(n267), .C1(n1657), .Y(n332) );
  CLKINVX1 U1445 ( .A(n286), .Y(n1001) );
  AOI222XL U1446 ( .A0(HI_mul[21]), .A1(n285), .B0(HI_div[21]), .B1(n273), 
        .C0(n260), .C1(n68), .Y(n286) );
  CLKINVX1 U1447 ( .A(n284), .Y(n1003) );
  AOI222XL U1448 ( .A0(HI_mul[20]), .A1(n285), .B0(HI_div[20]), .B1(n273), 
        .C0(n263), .C1(n69), .Y(n284) );
  CLKINVX1 U1449 ( .A(n280), .Y(n1007) );
  AOI222XL U1450 ( .A0(HI_mul[19]), .A1(n285), .B0(HI_div[19]), .B1(n277), 
        .C0(n265), .C1(n1683), .Y(n280) );
  CLKINVX1 U1451 ( .A(n278), .Y(n1009) );
  AOI222XL U1452 ( .A0(HI_mul[18]), .A1(n285), .B0(HI_div[18]), .B1(n275), 
        .C0(n265), .C1(n1682), .Y(n278) );
  CLKINVX1 U1453 ( .A(n276), .Y(n1011) );
  AOI222XL U1454 ( .A0(HI_mul[17]), .A1(n285), .B0(HI_div[17]), .B1(n273), 
        .C0(n265), .C1(n1681), .Y(n276) );
  CLKINVX1 U1455 ( .A(n274), .Y(n1013) );
  AOI222XL U1456 ( .A0(HI_mul[16]), .A1(n285), .B0(HI_div[16]), .B1(n277), 
        .C0(n265), .C1(n1680), .Y(n274) );
  CLKINVX1 U1457 ( .A(n272), .Y(n1015) );
  AOI222XL U1458 ( .A0(HI_mul[15]), .A1(n285), .B0(HI_div[15]), .B1(n275), 
        .C0(n265), .C1(n1679), .Y(n272) );
  CLKINVX1 U1459 ( .A(n270), .Y(n1282) );
  AOI222XL U1460 ( .A0(HI_mul[14]), .A1(n285), .B0(HI_div[14]), .B1(n271), 
        .C0(n265), .C1(n1678), .Y(n270) );
  CLKINVX1 U1461 ( .A(n268), .Y(n1283) );
  AOI222XL U1462 ( .A0(HI_mul[13]), .A1(n285), .B0(HI_div[13]), .B1(n271), 
        .C0(n265), .C1(n1677), .Y(n268) );
  CLKINVX1 U1463 ( .A(n266), .Y(n1284) );
  AOI222XL U1464 ( .A0(HI_mul[12]), .A1(n285), .B0(HI_div[12]), .B1(n271), 
        .C0(n265), .C1(n1676), .Y(n266) );
  CLKINVX1 U1465 ( .A(n382), .Y(n923) );
  AOI222XL U1466 ( .A0(LO_mul[7]), .A1(n279), .B0(LO_div[7]), .B1(n271), .C0(
        n267), .C1(n1651), .Y(n382) );
  CLKINVX1 U1467 ( .A(n380), .Y(n924) );
  AOI222XL U1468 ( .A0(LO_mul[6]), .A1(n279), .B0(LO_div[6]), .B1(n277), .C0(
        n269), .C1(n1650), .Y(n380) );
  CLKINVX1 U1469 ( .A(n264), .Y(n1285) );
  AOI222XL U1470 ( .A0(HI_mul[11]), .A1(n285), .B0(HI_div[11]), .B1(n259), 
        .C0(n265), .C1(n1675), .Y(n264) );
  CLKINVX1 U1471 ( .A(n262), .Y(n1286) );
  AOI222XL U1472 ( .A0(HI_mul[10]), .A1(n283), .B0(HI_div[10]), .B1(n273), 
        .C0(n265), .C1(n1674), .Y(n262) );
  CLKINVX1 U1473 ( .A(n322), .Y(n965) );
  AOI222XL U1474 ( .A0(HI_mul[9]), .A1(n283), .B0(HI_div[9]), .B1(n271), .C0(
        n265), .C1(n1673), .Y(n322) );
  CLKINVX1 U1475 ( .A(n320), .Y(n967) );
  AOI222XL U1476 ( .A0(HI_mul[8]), .A1(n283), .B0(HI_div[8]), .B1(n271), .C0(
        n267), .C1(n1672), .Y(n320) );
  CLKINVX1 U1477 ( .A(n330), .Y(n957) );
  AOI222XL U1478 ( .A0(LO_mul[12]), .A1(n281), .B0(LO_div[12]), .B1(n271), 
        .C0(n269), .C1(n1656), .Y(n330) );
  CLKINVX1 U1479 ( .A(n328), .Y(n959) );
  AOI222XL U1480 ( .A0(LO_mul[11]), .A1(n281), .B0(LO_div[11]), .B1(n259), 
        .C0(n269), .C1(n1655), .Y(n328) );
  CLKINVX1 U1481 ( .A(take), .Y(n1470) );
  CLKINVX1 U1482 ( .A(n318), .Y(n969) );
  AOI222XL U1483 ( .A0(HI_mul[7]), .A1(n283), .B0(HI_div[7]), .B1(n271), .C0(
        n263), .C1(n1671), .Y(n318) );
  CLKINVX1 U1484 ( .A(n316), .Y(n971) );
  AOI222XL U1485 ( .A0(HI_mul[6]), .A1(n283), .B0(HI_div[6]), .B1(n271), .C0(
        n263), .C1(n1670), .Y(n316) );
  CLKINVX1 U1486 ( .A(n314), .Y(n973) );
  AOI222XL U1487 ( .A0(HI_mul[5]), .A1(n283), .B0(HI_div[5]), .B1(n271), .C0(
        n263), .C1(n1669), .Y(n314) );
  CLKINVX1 U1488 ( .A(n312), .Y(n975) );
  AOI222XL U1489 ( .A0(HI_mul[4]), .A1(n283), .B0(HI_div[4]), .B1(n271), .C0(
        n263), .C1(n1668), .Y(n312) );
  CLKINVX1 U1490 ( .A(n310), .Y(n977) );
  AOI222XL U1491 ( .A0(HI_mul[3]), .A1(n283), .B0(HI_div[3]), .B1(n271), .C0(
        n269), .C1(n1667), .Y(n310) );
  CLKINVX1 U1492 ( .A(n304), .Y(n983) );
  AOI222XL U1493 ( .A0(HI_mul[2]), .A1(n283), .B0(HI_div[2]), .B1(n273), .C0(
        n263), .C1(n1666), .Y(n304) );
  CLKINVX1 U1494 ( .A(n282), .Y(n1005) );
  AOI222XL U1495 ( .A0(HI_mul[1]), .A1(n285), .B0(HI_div[1]), .B1(n259), .C0(
        n265), .C1(n1665), .Y(n282) );
  CLKINVX1 U1496 ( .A(n257), .Y(n1287) );
  AOI222XL U1497 ( .A0(HI_mul[0]), .A1(n281), .B0(HI_div[0]), .B1(n273), .C0(
        n265), .C1(n1664), .Y(n257) );
  CLKINVX1 U1498 ( .A(n326), .Y(n961) );
  AOI222XL U1499 ( .A0(LO_mul[10]), .A1(n283), .B0(LO_div[10]), .B1(n271), 
        .C0(n265), .C1(n1654), .Y(n326) );
  CLKINVX1 U1500 ( .A(n386), .Y(n921) );
  AOI222XL U1501 ( .A0(LO_mul[9]), .A1(n279), .B0(LO_div[9]), .B1(n275), .C0(
        n263), .C1(n1653), .Y(n386) );
  CLKINVX1 U1502 ( .A(n384), .Y(n922) );
  AOI222XL U1503 ( .A0(LO_mul[8]), .A1(n279), .B0(LO_div[8]), .B1(n271), .C0(
        n263), .C1(n1652), .Y(n384) );
  CLKINVX1 U1504 ( .A(n378), .Y(n925) );
  AOI222XL U1505 ( .A0(LO_mul[5]), .A1(n279), .B0(LO_div[5]), .B1(n277), .C0(
        n269), .C1(n1649), .Y(n378) );
  CLKINVX1 U1506 ( .A(n376), .Y(n926) );
  AOI222XL U1507 ( .A0(LO_mul[4]), .A1(n279), .B0(LO_div[4]), .B1(n277), .C0(
        n269), .C1(n1648), .Y(n376) );
  CLKINVX1 U1508 ( .A(n374), .Y(n927) );
  AOI222XL U1509 ( .A0(LO_mul[3]), .A1(n279), .B0(LO_div[3]), .B1(n277), .C0(
        n269), .C1(n1647), .Y(n374) );
  CLKINVX1 U1510 ( .A(n368), .Y(n930) );
  AOI222XL U1511 ( .A0(LO_mul[2]), .A1(n279), .B0(LO_div[2]), .B1(n277), .C0(
        n269), .C1(n1646), .Y(n368) );
  CLKINVX1 U1512 ( .A(n346), .Y(n941) );
  AOI222XL U1513 ( .A0(LO_mul[1]), .A1(n281), .B0(LO_div[1]), .B1(n275), .C0(
        n267), .C1(n1645), .Y(n346) );
  CLKINVX1 U1514 ( .A(n324), .Y(n963) );
  AOI222XL U1515 ( .A0(LO_mul[0]), .A1(n283), .B0(LO_div[0]), .B1(n271), .C0(
        n269), .C1(n1644), .Y(n324) );
  CLKBUFX3 U1516 ( .A(n259), .Y(n271) );
  NOR3X1 U1517 ( .A(n1397), .B(stall_div), .C(n279), .Y(n259) );
endmodule


module cache_0 ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   proc_addr_1, proc_addr_0, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         \tag_r[7][18] , \tag_r[7][17] , \tag_r[7][15] , \tag_r[7][14] ,
         \tag_r[7][13] , \tag_r[7][12] , \tag_r[7][11] , \tag_r[7][6] ,
         \tag_r[7][4] , \tag_r[7][3] , \tag_r[7][2] , \tag_r[7][1] ,
         \tag_r[7][0] , \tag_r[6][18] , \tag_r[6][17] , \tag_r[6][16] ,
         \tag_r[6][15] , \tag_r[6][14] , \tag_r[6][13] , \tag_r[6][12] ,
         \tag_r[6][6] , \tag_r[6][4] , \tag_r[6][3] , \tag_r[6][2] ,
         \tag_r[6][1] , \tag_r[6][0] , \tag_r[5][18] , \tag_r[5][17] ,
         \tag_r[5][16] , \tag_r[5][15] , \tag_r[5][14] , \tag_r[5][13] ,
         \tag_r[5][12] , \tag_r[5][6] , \tag_r[5][4] , \tag_r[5][3] ,
         \tag_r[5][2] , \tag_r[5][1] , \tag_r[5][0] , \tag_r[4][18] ,
         \tag_r[4][17] , \tag_r[4][16] , \tag_r[4][15] , \tag_r[4][14] ,
         \tag_r[4][13] , \tag_r[4][12] , \tag_r[4][6] , \tag_r[4][4] ,
         \tag_r[4][3] , \tag_r[4][2] , \tag_r[4][1] , \tag_r[4][0] ,
         \tag_r[3][18] , \tag_r[3][17] , \tag_r[3][16] , \tag_r[3][15] ,
         \tag_r[3][14] , \tag_r[3][13] , \tag_r[3][12] , \tag_r[3][6] ,
         \tag_r[3][4] , \tag_r[3][3] , \tag_r[3][2] , \tag_r[3][1] ,
         \tag_r[3][0] , \tag_r[2][18] , \tag_r[2][17] , \tag_r[2][16] ,
         \tag_r[2][15] , \tag_r[2][14] , \tag_r[2][13] , \tag_r[2][12] ,
         \tag_r[2][6] , \tag_r[2][4] , \tag_r[2][3] , \tag_r[2][2] ,
         \tag_r[2][1] , \tag_r[2][0] , \tag_r[1][18] , \tag_r[1][17] ,
         \tag_r[1][16] , \tag_r[1][15] , \tag_r[1][14] , \tag_r[1][13] ,
         \tag_r[1][12] , \tag_r[1][6] , \tag_r[1][4] , \tag_r[1][3] ,
         \tag_r[1][2] , \tag_r[1][1] , \tag_r[1][0] , \tag_r[0][18] ,
         \tag_r[0][17] , \tag_r[0][15] , \tag_r[0][14] , \tag_r[0][13] ,
         \tag_r[0][12] , \tag_r[0][11] , \tag_r[0][6] , \tag_r[0][4] ,
         \tag_r[0][3] , \tag_r[0][2] , \tag_r[0][1] , \tag_r[0][0] ,
         \state_r[0] , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n61, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1360, n1361, n1362,
         n1364, n1366, n1367, n1368, n1369, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1547,
         n1548, n1549, n1551, n1553, n1554, n1555, n1556, n1557, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1694, n1698, n1699, n1700, n1702, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1363, n1365, n1370, n1528, n1546,
         n1550, n1552, n1558, n1580, n1693, n1695, n1696, n1697, n1701, n1703,
         n1704, n2628, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418;
  assign proc_addr_1 = proc_addr[1];
  assign proc_addr_0 = proc_addr[0];

  DFFRX1 \block_r_reg[1][9]  ( .D(n3639), .CK(clk), .RN(n4285), .QN(n951) );
  DFFRX1 \block_r_reg[1][8]  ( .D(n3640), .CK(clk), .RN(n4284), .QN(n952) );
  DFFRX1 \block_r_reg[1][7]  ( .D(n3641), .CK(clk), .RN(n4284), .QN(n953) );
  DFFRX1 \block_r_reg[1][6]  ( .D(n3642), .CK(clk), .RN(n4283), .QN(n954) );
  DFFRX1 \block_r_reg[5][5]  ( .D(n3131), .CK(clk), .RN(n4283), .QN(n443) );
  DFFRX1 \block_r_reg[1][5]  ( .D(n3643), .CK(clk), .RN(n4282), .QN(n955) );
  DFFRX1 \block_r_reg[5][4]  ( .D(n3132), .CK(clk), .RN(n4282), .QN(n444) );
  DFFRX1 \block_r_reg[1][4]  ( .D(n3644), .CK(clk), .RN(n4282), .QN(n956) );
  DFFRX1 \block_r_reg[5][3]  ( .D(n3133), .CK(clk), .RN(n4281), .QN(n445) );
  DFFRX1 \block_r_reg[1][3]  ( .D(n3645), .CK(clk), .RN(n4281), .QN(n957) );
  DFFRX1 \block_r_reg[5][2]  ( .D(n3134), .CK(clk), .RN(n4281), .QN(n446) );
  DFFRX1 \block_r_reg[1][2]  ( .D(n3646), .CK(clk), .RN(n4280), .QN(n958) );
  DFFRX1 \block_r_reg[5][1]  ( .D(n3135), .CK(clk), .RN(n4280), .QN(n447) );
  DFFRX1 \block_r_reg[1][1]  ( .D(n3647), .CK(clk), .RN(n4280), .QN(n959) );
  DFFRX1 \block_r_reg[5][0]  ( .D(n3136), .CK(clk), .RN(n4279), .QN(n448) );
  DFFRX1 \block_r_reg[1][0]  ( .D(n3648), .CK(clk), .RN(n4279), .QN(n960) );
  DFFRX1 \block_r_reg[1][127]  ( .D(n3521), .CK(clk), .RN(n4278), .QN(n833) );
  DFFRX1 \block_r_reg[1][126]  ( .D(n3522), .CK(clk), .RN(n4278), .QN(n834) );
  DFFRX1 \block_r_reg[1][125]  ( .D(n3523), .CK(clk), .RN(n4277), .QN(n835) );
  DFFRX1 \block_r_reg[1][124]  ( .D(n3524), .CK(clk), .RN(n4276), .QN(n836) );
  DFFRX1 \block_r_reg[1][123]  ( .D(n3525), .CK(clk), .RN(n4276), .QN(n837) );
  DFFRX1 \block_r_reg[1][122]  ( .D(n3526), .CK(clk), .RN(n4275), .QN(n838) );
  DFFRX1 \block_r_reg[1][121]  ( .D(n3527), .CK(clk), .RN(n4274), .QN(n839) );
  DFFRX1 \block_r_reg[1][120]  ( .D(n3528), .CK(clk), .RN(n4274), .QN(n840) );
  DFFRX1 \block_r_reg[1][119]  ( .D(n3529), .CK(clk), .RN(n4273), .QN(n841) );
  DFFRX1 \block_r_reg[1][118]  ( .D(n3530), .CK(clk), .RN(n4272), .QN(n842) );
  DFFRX1 \block_r_reg[1][117]  ( .D(n3531), .CK(clk), .RN(n4272), .QN(n843) );
  DFFRX1 \block_r_reg[1][116]  ( .D(n3532), .CK(clk), .RN(n4271), .QN(n844) );
  DFFRX1 \block_r_reg[1][115]  ( .D(n3533), .CK(clk), .RN(n4270), .QN(n845) );
  DFFRX1 \block_r_reg[1][114]  ( .D(n3534), .CK(clk), .RN(n4270), .QN(n846) );
  DFFRX1 \block_r_reg[1][113]  ( .D(n3535), .CK(clk), .RN(n4269), .QN(n847) );
  DFFRX1 \block_r_reg[1][112]  ( .D(n3536), .CK(clk), .RN(n4268), .QN(n848) );
  DFFRX1 \block_r_reg[1][111]  ( .D(n3537), .CK(clk), .RN(n4268), .QN(n849) );
  DFFRX1 \block_r_reg[1][110]  ( .D(n3538), .CK(clk), .RN(n4267), .QN(n850) );
  DFFRX1 \block_r_reg[1][109]  ( .D(n3539), .CK(clk), .RN(n4266), .QN(n851) );
  DFFRX1 \block_r_reg[1][108]  ( .D(n3540), .CK(clk), .RN(n4266), .QN(n852) );
  DFFRX1 \block_r_reg[1][107]  ( .D(n3541), .CK(clk), .RN(n4265), .QN(n853) );
  DFFRX1 \block_r_reg[1][106]  ( .D(n3542), .CK(clk), .RN(n4264), .QN(n854) );
  DFFRX1 \block_r_reg[1][105]  ( .D(n3543), .CK(clk), .RN(n4264), .QN(n855) );
  DFFRX1 \block_r_reg[5][104]  ( .D(n3032), .CK(clk), .RN(n4263), .QN(n344) );
  DFFRX1 \block_r_reg[1][104]  ( .D(n3544), .CK(clk), .RN(n4263), .QN(n856) );
  DFFRX1 \block_r_reg[5][103]  ( .D(n3033), .CK(clk), .RN(n4263), .QN(n345) );
  DFFRX1 \block_r_reg[1][103]  ( .D(n3545), .CK(clk), .RN(n4262), .QN(n857) );
  DFFRX1 \block_r_reg[5][102]  ( .D(n3034), .CK(clk), .RN(n4262), .QN(n346) );
  DFFRX1 \block_r_reg[1][102]  ( .D(n3546), .CK(clk), .RN(n4262), .QN(n858) );
  DFFRX1 \block_r_reg[5][101]  ( .D(n3035), .CK(clk), .RN(n4261), .QN(n347) );
  DFFRX1 \block_r_reg[1][101]  ( .D(n3547), .CK(clk), .RN(n4261), .QN(n859) );
  DFFRX1 \block_r_reg[5][100]  ( .D(n3036), .CK(clk), .RN(n4261), .QN(n348) );
  DFFRX1 \block_r_reg[1][100]  ( .D(n3548), .CK(clk), .RN(n4260), .QN(n860) );
  DFFRX1 \block_r_reg[5][99]  ( .D(n3037), .CK(clk), .RN(n4260), .QN(n349) );
  DFFRX1 \block_r_reg[1][99]  ( .D(n3549), .CK(clk), .RN(n4260), .QN(n861) );
  DFFRX1 \block_r_reg[5][98]  ( .D(n3038), .CK(clk), .RN(n4259), .QN(n350) );
  DFFRX1 \block_r_reg[1][98]  ( .D(n3550), .CK(clk), .RN(n4259), .QN(n862) );
  DFFRX1 \block_r_reg[5][97]  ( .D(n3039), .CK(clk), .RN(n4259), .QN(n351) );
  DFFRX1 \block_r_reg[1][97]  ( .D(n3551), .CK(clk), .RN(n4258), .QN(n863) );
  DFFRX1 \block_r_reg[5][96]  ( .D(n3040), .CK(clk), .RN(n4258), .QN(n352) );
  DFFRX1 \block_r_reg[1][96]  ( .D(n3552), .CK(clk), .RN(n4258), .QN(n864) );
  DFFRX1 \block_r_reg[5][95]  ( .D(n3041), .CK(clk), .RN(n4257), .QN(n353) );
  DFFRX1 \block_r_reg[1][95]  ( .D(n3553), .CK(clk), .RN(n4257), .QN(n865) );
  DFFRX1 \block_r_reg[5][94]  ( .D(n3042), .CK(clk), .RN(n4257), .QN(n354) );
  DFFRX1 \block_r_reg[1][94]  ( .D(n3554), .CK(clk), .RN(n4256), .QN(n866) );
  DFFRX1 \block_r_reg[5][93]  ( .D(n3043), .CK(clk), .RN(n4256), .QN(n355) );
  DFFRX1 \block_r_reg[1][93]  ( .D(n3555), .CK(clk), .RN(n4256), .QN(n867) );
  DFFRX1 \block_r_reg[5][92]  ( .D(n3044), .CK(clk), .RN(n4255), .QN(n356) );
  DFFRX1 \block_r_reg[1][92]  ( .D(n3556), .CK(clk), .RN(n4255), .QN(n868) );
  DFFRX1 \block_r_reg[5][91]  ( .D(n3045), .CK(clk), .RN(n4255), .QN(n357) );
  DFFRX1 \block_r_reg[1][91]  ( .D(n3557), .CK(clk), .RN(n4254), .QN(n869) );
  DFFRX1 \block_r_reg[5][90]  ( .D(n3046), .CK(clk), .RN(n4254), .QN(n358) );
  DFFRX1 \block_r_reg[1][90]  ( .D(n3558), .CK(clk), .RN(n4254), .QN(n870) );
  DFFRX1 \block_r_reg[5][89]  ( .D(n3047), .CK(clk), .RN(n4253), .QN(n359) );
  DFFRX1 \block_r_reg[1][89]  ( .D(n3559), .CK(clk), .RN(n4253), .QN(n871) );
  DFFRX1 \block_r_reg[1][88]  ( .D(n3560), .CK(clk), .RN(n4252), .QN(n872) );
  DFFRX1 \block_r_reg[1][87]  ( .D(n3561), .CK(clk), .RN(n4252), .QN(n873) );
  DFFRX1 \block_r_reg[1][86]  ( .D(n3562), .CK(clk), .RN(n4251), .QN(n874) );
  DFFRX1 \block_r_reg[1][85]  ( .D(n3563), .CK(clk), .RN(n4250), .QN(n875) );
  DFFRX1 \block_r_reg[1][84]  ( .D(n3564), .CK(clk), .RN(n4250), .QN(n876) );
  DFFRX1 \block_r_reg[1][83]  ( .D(n3565), .CK(clk), .RN(n4249), .QN(n877) );
  DFFRX1 \block_r_reg[1][82]  ( .D(n3566), .CK(clk), .RN(n4248), .QN(n878) );
  DFFRX1 \block_r_reg[1][81]  ( .D(n3567), .CK(clk), .RN(n4248), .QN(n879) );
  DFFRX1 \block_r_reg[1][80]  ( .D(n3568), .CK(clk), .RN(n4247), .QN(n880) );
  DFFRX1 \block_r_reg[1][79]  ( .D(n3569), .CK(clk), .RN(n4246), .QN(n881) );
  DFFRX1 \block_r_reg[1][78]  ( .D(n3570), .CK(clk), .RN(n4246), .QN(n882) );
  DFFRX1 \block_r_reg[1][77]  ( .D(n3571), .CK(clk), .RN(n4245), .QN(n883) );
  DFFRX1 \block_r_reg[1][76]  ( .D(n3572), .CK(clk), .RN(n4244), .QN(n884) );
  DFFRX1 \block_r_reg[1][75]  ( .D(n3573), .CK(clk), .RN(n4244), .QN(n885) );
  DFFRX1 \block_r_reg[1][74]  ( .D(n3574), .CK(clk), .RN(n4243), .QN(n886) );
  DFFRX1 \block_r_reg[1][73]  ( .D(n3575), .CK(clk), .RN(n4242), .QN(n887) );
  DFFRX1 \block_r_reg[1][72]  ( .D(n3576), .CK(clk), .RN(n4242), .QN(n888) );
  DFFRX1 \block_r_reg[1][71]  ( .D(n3577), .CK(clk), .RN(n4241), .QN(n889) );
  DFFRX1 \block_r_reg[1][70]  ( .D(n3578), .CK(clk), .RN(n4240), .QN(n890) );
  DFFRX1 \block_r_reg[1][69]  ( .D(n3579), .CK(clk), .RN(n4240), .QN(n891) );
  DFFRX1 \block_r_reg[1][68]  ( .D(n3580), .CK(clk), .RN(n4239), .QN(n892) );
  DFFRX1 \block_r_reg[1][67]  ( .D(n3581), .CK(clk), .RN(n4238), .QN(n893) );
  DFFRX1 \block_r_reg[1][66]  ( .D(n3582), .CK(clk), .RN(n4238), .QN(n894) );
  DFFRX1 \block_r_reg[1][65]  ( .D(n3583), .CK(clk), .RN(n4237), .QN(n895) );
  DFFRX1 \block_r_reg[1][64]  ( .D(n3584), .CK(clk), .RN(n4236), .QN(n896) );
  DFFRX1 \block_r_reg[1][63]  ( .D(n3585), .CK(clk), .RN(n4236), .QN(n897) );
  DFFRX1 \block_r_reg[1][62]  ( .D(n3586), .CK(clk), .RN(n4235), .QN(n898) );
  DFFRX1 \block_r_reg[1][61]  ( .D(n3587), .CK(clk), .RN(n4234), .QN(n899) );
  DFFRX1 \block_r_reg[1][60]  ( .D(n3588), .CK(clk), .RN(n4234), .QN(n900) );
  DFFRX1 \block_r_reg[1][59]  ( .D(n3589), .CK(clk), .RN(n4233), .QN(n901) );
  DFFRX1 \block_r_reg[1][58]  ( .D(n3590), .CK(clk), .RN(n4232), .QN(n902) );
  DFFRX1 \block_r_reg[1][57]  ( .D(n3591), .CK(clk), .RN(n4232), .QN(n903) );
  DFFRX1 \block_r_reg[1][56]  ( .D(n3592), .CK(clk), .RN(n4231), .QN(n904) );
  DFFRX1 \block_r_reg[1][55]  ( .D(n3593), .CK(clk), .RN(n4230), .QN(n905) );
  DFFRX1 \block_r_reg[1][54]  ( .D(n3594), .CK(clk), .RN(n4230), .QN(n906) );
  DFFRX1 \block_r_reg[1][53]  ( .D(n3595), .CK(clk), .RN(n4229), .QN(n907) );
  DFFRX1 \block_r_reg[1][52]  ( .D(n3596), .CK(clk), .RN(n4228), .QN(n908) );
  DFFRX1 \block_r_reg[1][51]  ( .D(n3597), .CK(clk), .RN(n4228), .QN(n909) );
  DFFRX1 \block_r_reg[1][50]  ( .D(n3598), .CK(clk), .RN(n4227), .QN(n910) );
  DFFRX1 \block_r_reg[1][49]  ( .D(n3599), .CK(clk), .RN(n4226), .QN(n911) );
  DFFRX1 \block_r_reg[1][48]  ( .D(n3600), .CK(clk), .RN(n4226), .QN(n912) );
  DFFRX1 \block_r_reg[1][47]  ( .D(n3601), .CK(clk), .RN(n4225), .QN(n913) );
  DFFRX1 \block_r_reg[1][46]  ( .D(n3602), .CK(clk), .RN(n4224), .QN(n914) );
  DFFRX1 \block_r_reg[1][45]  ( .D(n3603), .CK(clk), .RN(n4224), .QN(n915) );
  DFFRX1 \block_r_reg[1][44]  ( .D(n3604), .CK(clk), .RN(n4223), .QN(n916) );
  DFFRX1 \block_r_reg[1][43]  ( .D(n3605), .CK(clk), .RN(n4222), .QN(n917) );
  DFFRX1 \block_r_reg[1][42]  ( .D(n3606), .CK(clk), .RN(n4222), .QN(n918) );
  DFFRX1 \block_r_reg[1][41]  ( .D(n3607), .CK(clk), .RN(n4221), .QN(n919) );
  DFFRX1 \block_r_reg[1][40]  ( .D(n3608), .CK(clk), .RN(n4220), .QN(n920) );
  DFFRX1 \block_r_reg[1][39]  ( .D(n3609), .CK(clk), .RN(n4220), .QN(n921) );
  DFFRX1 \block_r_reg[1][38]  ( .D(n3610), .CK(clk), .RN(n4219), .QN(n922) );
  DFFRX1 \block_r_reg[1][37]  ( .D(n3611), .CK(clk), .RN(n4218), .QN(n923) );
  DFFRX1 \block_r_reg[1][36]  ( .D(n3612), .CK(clk), .RN(n4218), .QN(n924) );
  DFFRX1 \block_r_reg[1][35]  ( .D(n3613), .CK(clk), .RN(n4217), .QN(n925) );
  DFFRX1 \block_r_reg[1][34]  ( .D(n3614), .CK(clk), .RN(n4216), .QN(n926) );
  DFFRX1 \block_r_reg[1][33]  ( .D(n3615), .CK(clk), .RN(n4216), .QN(n927) );
  DFFRX1 \block_r_reg[1][32]  ( .D(n3616), .CK(clk), .RN(n4215), .QN(n928) );
  DFFRX1 \block_r_reg[1][31]  ( .D(n3617), .CK(clk), .RN(n4214), .QN(n929) );
  DFFRX1 \block_r_reg[1][30]  ( .D(n3618), .CK(clk), .RN(n4214), .QN(n930) );
  DFFRX1 \block_r_reg[1][29]  ( .D(n3619), .CK(clk), .RN(n4213), .QN(n931) );
  DFFRX1 \block_r_reg[1][28]  ( .D(n3620), .CK(clk), .RN(n4212), .QN(n932) );
  DFFRX1 \block_r_reg[1][27]  ( .D(n3621), .CK(clk), .RN(n4212), .QN(n933) );
  DFFRX1 \block_r_reg[1][26]  ( .D(n3622), .CK(clk), .RN(n4211), .QN(n934) );
  DFFRX1 \block_r_reg[1][25]  ( .D(n3623), .CK(clk), .RN(n4210), .QN(n935) );
  DFFRX1 \block_r_reg[1][24]  ( .D(n3624), .CK(clk), .RN(n4210), .QN(n936) );
  DFFRX1 \block_r_reg[1][23]  ( .D(n3625), .CK(clk), .RN(n4209), .QN(n937) );
  DFFRX1 \block_r_reg[1][22]  ( .D(n3626), .CK(clk), .RN(n4208), .QN(n938) );
  DFFRX1 \block_r_reg[1][21]  ( .D(n3627), .CK(clk), .RN(n4208), .QN(n939) );
  DFFRX1 \block_r_reg[1][20]  ( .D(n3628), .CK(clk), .RN(n4207), .QN(n940) );
  DFFRX1 \block_r_reg[1][19]  ( .D(n3629), .CK(clk), .RN(n4206), .QN(n941) );
  DFFRX1 \block_r_reg[1][18]  ( .D(n3630), .CK(clk), .RN(n4206), .QN(n942) );
  DFFRX1 \block_r_reg[7][17]  ( .D(n2863), .CK(clk), .RN(n4291), .QN(n175) );
  DFFRX1 \block_r_reg[5][17]  ( .D(n3119), .CK(clk), .RN(n4291), .QN(n431) );
  DFFRX1 \block_r_reg[3][17]  ( .D(n3375), .CK(clk), .RN(n4290), .QN(n687) );
  DFFRX1 \block_r_reg[7][16]  ( .D(n2864), .CK(clk), .RN(n4290), .QN(n176) );
  DFFRX1 \block_r_reg[5][16]  ( .D(n3120), .CK(clk), .RN(n4290), .QN(n432) );
  DFFRX1 \block_r_reg[3][16]  ( .D(n3376), .CK(clk), .RN(n4290), .QN(n688) );
  DFFRX1 \block_r_reg[7][15]  ( .D(n2865), .CK(clk), .RN(n4289), .QN(n177) );
  DFFRX1 \block_r_reg[5][15]  ( .D(n3121), .CK(clk), .RN(n4289), .QN(n433) );
  DFFRX1 \block_r_reg[3][15]  ( .D(n3377), .CK(clk), .RN(n4289), .QN(n689) );
  DFFRX1 \block_r_reg[7][14]  ( .D(n2866), .CK(clk), .RN(n4289), .QN(n178) );
  DFFRX1 \block_r_reg[5][14]  ( .D(n3122), .CK(clk), .RN(n4289), .QN(n434) );
  DFFRX1 \block_r_reg[3][14]  ( .D(n3378), .CK(clk), .RN(n4288), .QN(n690) );
  DFFRX1 \block_r_reg[7][13]  ( .D(n2867), .CK(clk), .RN(n4288), .QN(n179) );
  DFFRX1 \block_r_reg[5][13]  ( .D(n3123), .CK(clk), .RN(n4288), .QN(n435) );
  DFFRX1 \block_r_reg[3][13]  ( .D(n3379), .CK(clk), .RN(n4288), .QN(n691) );
  DFFRX1 \block_r_reg[7][12]  ( .D(n2868), .CK(clk), .RN(n4287), .QN(n180) );
  DFFRX1 \block_r_reg[5][12]  ( .D(n3124), .CK(clk), .RN(n4287), .QN(n436) );
  DFFRX1 \block_r_reg[3][12]  ( .D(n3380), .CK(clk), .RN(n4287), .QN(n692) );
  DFFRX1 \block_r_reg[7][11]  ( .D(n2869), .CK(clk), .RN(n4287), .QN(n181) );
  DFFRX1 \block_r_reg[5][11]  ( .D(n3125), .CK(clk), .RN(n4287), .QN(n437) );
  DFFRX1 \block_r_reg[3][11]  ( .D(n3381), .CK(clk), .RN(n4286), .QN(n693) );
  DFFRX1 \block_r_reg[7][10]  ( .D(n2870), .CK(clk), .RN(n4286), .QN(n182) );
  DFFRX1 \block_r_reg[5][10]  ( .D(n3126), .CK(clk), .RN(n4286), .QN(n438) );
  DFFRX1 \block_r_reg[3][10]  ( .D(n3382), .CK(clk), .RN(n4286), .QN(n694) );
  DFFRX1 \block_r_reg[7][9]  ( .D(n2871), .CK(clk), .RN(n4285), .QN(n183) );
  DFFRX1 \block_r_reg[5][9]  ( .D(n3127), .CK(clk), .RN(n4285), .QN(n439) );
  DFFRX1 \block_r_reg[3][9]  ( .D(n3383), .CK(clk), .RN(n4285), .QN(n695) );
  DFFRX1 \block_r_reg[7][8]  ( .D(n2872), .CK(clk), .RN(n4285), .QN(n184) );
  DFFRX1 \block_r_reg[5][8]  ( .D(n3128), .CK(clk), .RN(n4285), .QN(n440) );
  DFFRX1 \block_r_reg[3][8]  ( .D(n3384), .CK(clk), .RN(n4284), .QN(n696) );
  DFFRX1 \block_r_reg[7][7]  ( .D(n2873), .CK(clk), .RN(n4284), .QN(n185) );
  DFFRX1 \block_r_reg[5][7]  ( .D(n3129), .CK(clk), .RN(n4284), .QN(n441) );
  DFFRX1 \block_r_reg[3][7]  ( .D(n3385), .CK(clk), .RN(n4284), .QN(n697) );
  DFFRX1 \block_r_reg[7][6]  ( .D(n2874), .CK(clk), .RN(n4283), .QN(n186) );
  DFFRX1 \block_r_reg[5][6]  ( .D(n3130), .CK(clk), .RN(n4283), .QN(n442) );
  DFFRX1 \block_r_reg[3][6]  ( .D(n3386), .CK(clk), .RN(n4283), .QN(n698) );
  DFFRX1 \block_r_reg[7][5]  ( .D(n2875), .CK(clk), .RN(n4283), .QN(n187) );
  DFFRX1 \block_r_reg[3][5]  ( .D(n3387), .CK(clk), .RN(n4282), .QN(n699) );
  DFFRX1 \block_r_reg[7][4]  ( .D(n2876), .CK(clk), .RN(n4282), .QN(n188) );
  DFFRX1 \block_r_reg[3][4]  ( .D(n3388), .CK(clk), .RN(n4282), .QN(n700) );
  DFFRX1 \block_r_reg[7][3]  ( .D(n2877), .CK(clk), .RN(n4281), .QN(n189) );
  DFFRX1 \block_r_reg[3][3]  ( .D(n3389), .CK(clk), .RN(n4281), .QN(n701) );
  DFFRX1 \block_r_reg[7][2]  ( .D(n2878), .CK(clk), .RN(n4281), .QN(n190) );
  DFFRX1 \block_r_reg[3][2]  ( .D(n3390), .CK(clk), .RN(n4280), .QN(n702) );
  DFFRX1 \block_r_reg[7][1]  ( .D(n2879), .CK(clk), .RN(n4280), .QN(n191) );
  DFFRX1 \block_r_reg[3][1]  ( .D(n3391), .CK(clk), .RN(n4280), .QN(n703) );
  DFFRX1 \block_r_reg[7][0]  ( .D(n2880), .CK(clk), .RN(n4279), .QN(n192) );
  DFFRX1 \block_r_reg[3][0]  ( .D(n3392), .CK(clk), .RN(n4279), .QN(n704) );
  DFFRX1 \block_r_reg[7][127]  ( .D(n2753), .CK(clk), .RN(n4279), .QN(n65) );
  DFFRX1 \block_r_reg[5][127]  ( .D(n3009), .CK(clk), .RN(n4279), .QN(n321) );
  DFFRX1 \block_r_reg[4][127]  ( .D(n3137), .CK(clk), .RN(n4278), .QN(n449) );
  DFFRX1 \block_r_reg[3][127]  ( .D(n3265), .CK(clk), .RN(n4278), .QN(n577) );
  DFFRX1 \block_r_reg[7][126]  ( .D(n2754), .CK(clk), .RN(n4278), .QN(n66) );
  DFFRX1 \block_r_reg[5][126]  ( .D(n3010), .CK(clk), .RN(n4278), .QN(n322) );
  DFFRX1 \block_r_reg[4][126]  ( .D(n3138), .CK(clk), .RN(n4278), .QN(n450) );
  DFFRX1 \block_r_reg[3][126]  ( .D(n3266), .CK(clk), .RN(n4278), .QN(n578) );
  DFFRX1 \block_r_reg[7][125]  ( .D(n2755), .CK(clk), .RN(n4277), .QN(n67) );
  DFFRX1 \block_r_reg[5][125]  ( .D(n3011), .CK(clk), .RN(n4277), .QN(n323) );
  DFFRX1 \block_r_reg[4][125]  ( .D(n3139), .CK(clk), .RN(n4277), .QN(n451) );
  DFFRX1 \block_r_reg[3][125]  ( .D(n3267), .CK(clk), .RN(n4277), .QN(n579) );
  DFFRX1 \block_r_reg[7][124]  ( .D(n2756), .CK(clk), .RN(n4277), .QN(n68) );
  DFFRX1 \block_r_reg[5][124]  ( .D(n3012), .CK(clk), .RN(n4277), .QN(n324) );
  DFFRX1 \block_r_reg[4][124]  ( .D(n3140), .CK(clk), .RN(n4276), .QN(n452) );
  DFFRX1 \block_r_reg[3][124]  ( .D(n3268), .CK(clk), .RN(n4276), .QN(n580) );
  DFFRX1 \block_r_reg[7][123]  ( .D(n2757), .CK(clk), .RN(n4276), .QN(n69) );
  DFFRX1 \block_r_reg[5][123]  ( .D(n3013), .CK(clk), .RN(n4276), .QN(n325) );
  DFFRX1 \block_r_reg[4][123]  ( .D(n3141), .CK(clk), .RN(n4276), .QN(n453) );
  DFFRX1 \block_r_reg[3][123]  ( .D(n3269), .CK(clk), .RN(n4276), .QN(n581) );
  DFFRX1 \block_r_reg[7][122]  ( .D(n2758), .CK(clk), .RN(n4275), .QN(n70) );
  DFFRX1 \block_r_reg[5][122]  ( .D(n3014), .CK(clk), .RN(n4275), .QN(n326) );
  DFFRX1 \block_r_reg[4][122]  ( .D(n3142), .CK(clk), .RN(n4275), .QN(n454) );
  DFFRX1 \block_r_reg[3][122]  ( .D(n3270), .CK(clk), .RN(n4275), .QN(n582) );
  DFFRX1 \block_r_reg[7][121]  ( .D(n2759), .CK(clk), .RN(n4275), .QN(n71) );
  DFFRX1 \block_r_reg[5][121]  ( .D(n3015), .CK(clk), .RN(n4275), .QN(n327) );
  DFFRX1 \block_r_reg[4][121]  ( .D(n3143), .CK(clk), .RN(n4274), .QN(n455) );
  DFFRX1 \block_r_reg[3][121]  ( .D(n3271), .CK(clk), .RN(n4274), .QN(n583) );
  DFFRX1 \block_r_reg[7][120]  ( .D(n2760), .CK(clk), .RN(n4274), .QN(n72) );
  DFFRX1 \block_r_reg[5][120]  ( .D(n3016), .CK(clk), .RN(n4274), .QN(n328) );
  DFFRX1 \block_r_reg[4][120]  ( .D(n3144), .CK(clk), .RN(n4274), .QN(n456) );
  DFFRX1 \block_r_reg[3][120]  ( .D(n3272), .CK(clk), .RN(n4274), .QN(n584) );
  DFFRX1 \block_r_reg[7][119]  ( .D(n2761), .CK(clk), .RN(n4273), .QN(n73) );
  DFFRX1 \block_r_reg[5][119]  ( .D(n3017), .CK(clk), .RN(n4273), .QN(n329) );
  DFFRX1 \block_r_reg[4][119]  ( .D(n3145), .CK(clk), .RN(n4273), .QN(n457) );
  DFFRX1 \block_r_reg[3][119]  ( .D(n3273), .CK(clk), .RN(n4273), .QN(n585) );
  DFFRX1 \block_r_reg[7][118]  ( .D(n2762), .CK(clk), .RN(n4273), .QN(n74) );
  DFFRX1 \block_r_reg[5][118]  ( .D(n3018), .CK(clk), .RN(n4273), .QN(n330) );
  DFFRX1 \block_r_reg[4][118]  ( .D(n3146), .CK(clk), .RN(n4272), .QN(n458) );
  DFFRX1 \block_r_reg[3][118]  ( .D(n3274), .CK(clk), .RN(n4272), .QN(n586) );
  DFFRX1 \block_r_reg[7][117]  ( .D(n2763), .CK(clk), .RN(n4272), .QN(n75) );
  DFFRX1 \block_r_reg[5][117]  ( .D(n3019), .CK(clk), .RN(n4272), .QN(n331) );
  DFFRX1 \block_r_reg[3][117]  ( .D(n3275), .CK(clk), .RN(n4272), .QN(n587) );
  DFFRX1 \block_r_reg[7][116]  ( .D(n2764), .CK(clk), .RN(n4271), .QN(n76) );
  DFFRX1 \block_r_reg[5][116]  ( .D(n3020), .CK(clk), .RN(n4271), .QN(n332) );
  DFFRX1 \block_r_reg[3][116]  ( .D(n3276), .CK(clk), .RN(n4271), .QN(n588) );
  DFFRX1 \block_r_reg[7][115]  ( .D(n2765), .CK(clk), .RN(n4271), .QN(n77) );
  DFFRX1 \block_r_reg[5][115]  ( .D(n3021), .CK(clk), .RN(n4271), .QN(n333) );
  DFFRX1 \block_r_reg[3][115]  ( .D(n3277), .CK(clk), .RN(n4270), .QN(n589) );
  DFFRX1 \block_r_reg[7][114]  ( .D(n2766), .CK(clk), .RN(n4270), .QN(n78) );
  DFFRX1 \block_r_reg[5][114]  ( .D(n3022), .CK(clk), .RN(n4270), .QN(n334) );
  DFFRX1 \block_r_reg[3][114]  ( .D(n3278), .CK(clk), .RN(n4270), .QN(n590) );
  DFFRX1 \block_r_reg[7][113]  ( .D(n2767), .CK(clk), .RN(n4269), .QN(n79) );
  DFFRX1 \block_r_reg[5][113]  ( .D(n3023), .CK(clk), .RN(n4269), .QN(n335) );
  DFFRX1 \block_r_reg[3][113]  ( .D(n3279), .CK(clk), .RN(n4269), .QN(n591) );
  DFFRX1 \block_r_reg[7][112]  ( .D(n2768), .CK(clk), .RN(n4269), .QN(n80) );
  DFFRX1 \block_r_reg[5][112]  ( .D(n3024), .CK(clk), .RN(n4269), .QN(n336) );
  DFFRX1 \block_r_reg[3][112]  ( .D(n3280), .CK(clk), .RN(n4268), .QN(n592) );
  DFFRX1 \block_r_reg[7][111]  ( .D(n2769), .CK(clk), .RN(n4268), .QN(n81) );
  DFFRX1 \block_r_reg[5][111]  ( .D(n3025), .CK(clk), .RN(n4268), .QN(n337) );
  DFFRX1 \block_r_reg[3][111]  ( .D(n3281), .CK(clk), .RN(n4268), .QN(n593) );
  DFFRX1 \block_r_reg[7][110]  ( .D(n2770), .CK(clk), .RN(n4267), .QN(n82) );
  DFFRX1 \block_r_reg[5][110]  ( .D(n3026), .CK(clk), .RN(n4267), .QN(n338) );
  DFFRX1 \block_r_reg[3][110]  ( .D(n3282), .CK(clk), .RN(n4267), .QN(n594) );
  DFFRX1 \block_r_reg[7][109]  ( .D(n2771), .CK(clk), .RN(n4267), .QN(n83) );
  DFFRX1 \block_r_reg[5][109]  ( .D(n3027), .CK(clk), .RN(n4267), .QN(n339) );
  DFFRX1 \block_r_reg[3][109]  ( .D(n3283), .CK(clk), .RN(n4266), .QN(n595) );
  DFFRX1 \block_r_reg[7][108]  ( .D(n2772), .CK(clk), .RN(n4266), .QN(n84) );
  DFFRX1 \block_r_reg[5][108]  ( .D(n3028), .CK(clk), .RN(n4266), .QN(n340) );
  DFFRX1 \block_r_reg[3][108]  ( .D(n3284), .CK(clk), .RN(n4266), .QN(n596) );
  DFFRX1 \block_r_reg[7][107]  ( .D(n2773), .CK(clk), .RN(n4265), .QN(n85) );
  DFFRX1 \block_r_reg[5][107]  ( .D(n3029), .CK(clk), .RN(n4265), .QN(n341) );
  DFFRX1 \block_r_reg[3][107]  ( .D(n3285), .CK(clk), .RN(n4265), .QN(n597) );
  DFFRX1 \block_r_reg[7][106]  ( .D(n2774), .CK(clk), .RN(n4265), .QN(n86) );
  DFFRX1 \block_r_reg[5][106]  ( .D(n3030), .CK(clk), .RN(n4265), .QN(n342) );
  DFFRX1 \block_r_reg[3][106]  ( .D(n3286), .CK(clk), .RN(n4264), .QN(n598) );
  DFFRX1 \block_r_reg[7][105]  ( .D(n2775), .CK(clk), .RN(n4264), .QN(n87) );
  DFFRX1 \block_r_reg[5][105]  ( .D(n3031), .CK(clk), .RN(n4264), .QN(n343) );
  DFFRX1 \block_r_reg[3][105]  ( .D(n3287), .CK(clk), .RN(n4264), .QN(n599) );
  DFFRX1 \block_r_reg[7][104]  ( .D(n2776), .CK(clk), .RN(n4263), .QN(n88) );
  DFFRX1 \block_r_reg[3][104]  ( .D(n3288), .CK(clk), .RN(n4263), .QN(n600) );
  DFFRX1 \block_r_reg[7][103]  ( .D(n2777), .CK(clk), .RN(n4263), .QN(n89) );
  DFFRX1 \block_r_reg[3][103]  ( .D(n3289), .CK(clk), .RN(n4262), .QN(n601) );
  DFFRX1 \block_r_reg[7][102]  ( .D(n2778), .CK(clk), .RN(n4262), .QN(n90) );
  DFFRX1 \block_r_reg[3][102]  ( .D(n3290), .CK(clk), .RN(n4262), .QN(n602) );
  DFFRX1 \block_r_reg[7][101]  ( .D(n2779), .CK(clk), .RN(n4261), .QN(n91) );
  DFFRX1 \block_r_reg[3][101]  ( .D(n3291), .CK(clk), .RN(n4261), .QN(n603) );
  DFFRX1 \block_r_reg[7][100]  ( .D(n2780), .CK(clk), .RN(n4261), .QN(n92) );
  DFFRX1 \block_r_reg[3][100]  ( .D(n3292), .CK(clk), .RN(n4260), .QN(n604) );
  DFFRX1 \block_r_reg[7][99]  ( .D(n2781), .CK(clk), .RN(n4260), .QN(n93) );
  DFFRX1 \block_r_reg[3][99]  ( .D(n3293), .CK(clk), .RN(n4260), .QN(n605) );
  DFFRX1 \block_r_reg[7][98]  ( .D(n2782), .CK(clk), .RN(n4259), .QN(n94) );
  DFFRX1 \block_r_reg[3][98]  ( .D(n3294), .CK(clk), .RN(n4259), .QN(n606) );
  DFFRX1 \block_r_reg[7][97]  ( .D(n2783), .CK(clk), .RN(n4259), .QN(n95) );
  DFFRX1 \block_r_reg[3][97]  ( .D(n3295), .CK(clk), .RN(n4258), .QN(n607) );
  DFFRX1 \block_r_reg[7][96]  ( .D(n2784), .CK(clk), .RN(n4258), .QN(n96) );
  DFFRX1 \block_r_reg[3][96]  ( .D(n3296), .CK(clk), .RN(n4258), .QN(n608) );
  DFFRX1 \block_r_reg[7][95]  ( .D(n2785), .CK(clk), .RN(n4257), .QN(n97) );
  DFFRX1 \block_r_reg[3][95]  ( .D(n3297), .CK(clk), .RN(n4257), .QN(n609) );
  DFFRX1 \block_r_reg[7][94]  ( .D(n2786), .CK(clk), .RN(n4257), .QN(n98) );
  DFFRX1 \block_r_reg[3][94]  ( .D(n3298), .CK(clk), .RN(n4256), .QN(n610) );
  DFFRX1 \block_r_reg[7][93]  ( .D(n2787), .CK(clk), .RN(n4256), .QN(n99) );
  DFFRX1 \block_r_reg[3][93]  ( .D(n3299), .CK(clk), .RN(n4256), .QN(n611) );
  DFFRX1 \block_r_reg[7][92]  ( .D(n2788), .CK(clk), .RN(n4255), .QN(n100) );
  DFFRX1 \block_r_reg[3][92]  ( .D(n3300), .CK(clk), .RN(n4255), .QN(n612) );
  DFFRX1 \block_r_reg[7][91]  ( .D(n2789), .CK(clk), .RN(n4255), .QN(n101) );
  DFFRX1 \block_r_reg[3][91]  ( .D(n3301), .CK(clk), .RN(n4254), .QN(n613) );
  DFFRX1 \block_r_reg[7][90]  ( .D(n2790), .CK(clk), .RN(n4254), .QN(n102) );
  DFFRX1 \block_r_reg[3][90]  ( .D(n3302), .CK(clk), .RN(n4254), .QN(n614) );
  DFFRX1 \block_r_reg[7][89]  ( .D(n2791), .CK(clk), .RN(n4253), .QN(n103) );
  DFFRX1 \block_r_reg[3][89]  ( .D(n3303), .CK(clk), .RN(n4253), .QN(n615) );
  DFFRX1 \block_r_reg[7][88]  ( .D(n2792), .CK(clk), .RN(n4253), .QN(n104) );
  DFFRX1 \block_r_reg[5][88]  ( .D(n3048), .CK(clk), .RN(n4253), .QN(n360) );
  DFFRX1 \block_r_reg[3][88]  ( .D(n3304), .CK(clk), .RN(n4252), .QN(n616) );
  DFFRX1 \block_r_reg[7][87]  ( .D(n2793), .CK(clk), .RN(n4252), .QN(n105) );
  DFFRX1 \block_r_reg[5][87]  ( .D(n3049), .CK(clk), .RN(n4252), .QN(n361) );
  DFFRX1 \block_r_reg[3][87]  ( .D(n3305), .CK(clk), .RN(n4252), .QN(n617) );
  DFFRX1 \block_r_reg[7][86]  ( .D(n2794), .CK(clk), .RN(n4251), .QN(n106) );
  DFFRX1 \block_r_reg[5][86]  ( .D(n3050), .CK(clk), .RN(n4251), .QN(n362) );
  DFFRX1 \block_r_reg[3][86]  ( .D(n3306), .CK(clk), .RN(n4251), .QN(n618) );
  DFFRX1 \block_r_reg[7][85]  ( .D(n2795), .CK(clk), .RN(n4251), .QN(n107) );
  DFFRX1 \block_r_reg[5][85]  ( .D(n3051), .CK(clk), .RN(n4251), .QN(n363) );
  DFFRX1 \block_r_reg[3][85]  ( .D(n3307), .CK(clk), .RN(n4250), .QN(n619) );
  DFFRX1 \block_r_reg[7][84]  ( .D(n2796), .CK(clk), .RN(n4250), .QN(n108) );
  DFFRX1 \block_r_reg[5][84]  ( .D(n3052), .CK(clk), .RN(n4250), .QN(n364) );
  DFFRX1 \block_r_reg[3][84]  ( .D(n3308), .CK(clk), .RN(n4250), .QN(n620) );
  DFFRX1 \block_r_reg[7][83]  ( .D(n2797), .CK(clk), .RN(n4249), .QN(n109) );
  DFFRX1 \block_r_reg[5][83]  ( .D(n3053), .CK(clk), .RN(n4249), .QN(n365) );
  DFFRX1 \block_r_reg[3][83]  ( .D(n3309), .CK(clk), .RN(n4249), .QN(n621) );
  DFFRX1 \block_r_reg[7][82]  ( .D(n2798), .CK(clk), .RN(n4249), .QN(n110) );
  DFFRX1 \block_r_reg[5][82]  ( .D(n3054), .CK(clk), .RN(n4249), .QN(n366) );
  DFFRX1 \block_r_reg[3][82]  ( .D(n3310), .CK(clk), .RN(n4248), .QN(n622) );
  DFFRX1 \block_r_reg[7][81]  ( .D(n2799), .CK(clk), .RN(n4248), .QN(n111) );
  DFFRX1 \block_r_reg[5][81]  ( .D(n3055), .CK(clk), .RN(n4248), .QN(n367) );
  DFFRX1 \block_r_reg[3][81]  ( .D(n3311), .CK(clk), .RN(n4248), .QN(n623) );
  DFFRX1 \block_r_reg[7][80]  ( .D(n2800), .CK(clk), .RN(n4247), .QN(n112) );
  DFFRX1 \block_r_reg[5][80]  ( .D(n3056), .CK(clk), .RN(n4247), .QN(n368) );
  DFFRX1 \block_r_reg[3][80]  ( .D(n3312), .CK(clk), .RN(n4247), .QN(n624) );
  DFFRX1 \block_r_reg[7][79]  ( .D(n2801), .CK(clk), .RN(n4247), .QN(n113) );
  DFFRX1 \block_r_reg[5][79]  ( .D(n3057), .CK(clk), .RN(n4247), .QN(n369) );
  DFFRX1 \block_r_reg[3][79]  ( .D(n3313), .CK(clk), .RN(n4246), .QN(n625) );
  DFFRX1 \block_r_reg[7][78]  ( .D(n2802), .CK(clk), .RN(n4246), .QN(n114) );
  DFFRX1 \block_r_reg[5][78]  ( .D(n3058), .CK(clk), .RN(n4246), .QN(n370) );
  DFFRX1 \block_r_reg[3][78]  ( .D(n3314), .CK(clk), .RN(n4246), .QN(n626) );
  DFFRX1 \block_r_reg[7][77]  ( .D(n2803), .CK(clk), .RN(n4245), .QN(n115) );
  DFFRX1 \block_r_reg[5][77]  ( .D(n3059), .CK(clk), .RN(n4245), .QN(n371) );
  DFFRX1 \block_r_reg[3][77]  ( .D(n3315), .CK(clk), .RN(n4245), .QN(n627) );
  DFFRX1 \block_r_reg[7][76]  ( .D(n2804), .CK(clk), .RN(n4245), .QN(n116) );
  DFFRX1 \block_r_reg[5][76]  ( .D(n3060), .CK(clk), .RN(n4245), .QN(n372) );
  DFFRX1 \block_r_reg[3][76]  ( .D(n3316), .CK(clk), .RN(n4244), .QN(n628) );
  DFFRX1 \block_r_reg[7][75]  ( .D(n2805), .CK(clk), .RN(n4244), .QN(n117) );
  DFFRX1 \block_r_reg[5][75]  ( .D(n3061), .CK(clk), .RN(n4244), .QN(n373) );
  DFFRX1 \block_r_reg[3][75]  ( .D(n3317), .CK(clk), .RN(n4244), .QN(n629) );
  DFFRX1 \block_r_reg[7][74]  ( .D(n2806), .CK(clk), .RN(n4243), .QN(n118) );
  DFFRX1 \block_r_reg[5][74]  ( .D(n3062), .CK(clk), .RN(n4243), .QN(n374) );
  DFFRX1 \block_r_reg[3][74]  ( .D(n3318), .CK(clk), .RN(n4243), .QN(n630) );
  DFFRX1 \block_r_reg[7][73]  ( .D(n2807), .CK(clk), .RN(n4243), .QN(n119) );
  DFFRX1 \block_r_reg[5][73]  ( .D(n3063), .CK(clk), .RN(n4243), .QN(n375) );
  DFFRX1 \block_r_reg[3][73]  ( .D(n3319), .CK(clk), .RN(n4242), .QN(n631) );
  DFFRX1 \block_r_reg[7][72]  ( .D(n2808), .CK(clk), .RN(n4242), .QN(n120) );
  DFFRX1 \block_r_reg[5][72]  ( .D(n3064), .CK(clk), .RN(n4242), .QN(n376) );
  DFFRX1 \block_r_reg[3][72]  ( .D(n3320), .CK(clk), .RN(n4242), .QN(n632) );
  DFFRX1 \block_r_reg[7][71]  ( .D(n2809), .CK(clk), .RN(n4241), .QN(n121) );
  DFFRX1 \block_r_reg[5][71]  ( .D(n3065), .CK(clk), .RN(n4241), .QN(n377) );
  DFFRX1 \block_r_reg[3][71]  ( .D(n3321), .CK(clk), .RN(n4241), .QN(n633) );
  DFFRX1 \block_r_reg[7][70]  ( .D(n2810), .CK(clk), .RN(n4241), .QN(n122) );
  DFFRX1 \block_r_reg[5][70]  ( .D(n3066), .CK(clk), .RN(n4241), .QN(n378) );
  DFFRX1 \block_r_reg[3][70]  ( .D(n3322), .CK(clk), .RN(n4240), .QN(n634) );
  DFFRX1 \block_r_reg[7][69]  ( .D(n2811), .CK(clk), .RN(n4240), .QN(n123) );
  DFFRX1 \block_r_reg[5][69]  ( .D(n3067), .CK(clk), .RN(n4240), .QN(n379) );
  DFFRX1 \block_r_reg[3][69]  ( .D(n3323), .CK(clk), .RN(n4240), .QN(n635) );
  DFFRX1 \block_r_reg[7][68]  ( .D(n2812), .CK(clk), .RN(n4239), .QN(n124) );
  DFFRX1 \block_r_reg[5][68]  ( .D(n3068), .CK(clk), .RN(n4239), .QN(n380) );
  DFFRX1 \block_r_reg[3][68]  ( .D(n3324), .CK(clk), .RN(n4239), .QN(n636) );
  DFFRX1 \block_r_reg[7][67]  ( .D(n2813), .CK(clk), .RN(n4239), .QN(n125) );
  DFFRX1 \block_r_reg[5][67]  ( .D(n3069), .CK(clk), .RN(n4239), .QN(n381) );
  DFFRX1 \block_r_reg[3][67]  ( .D(n3325), .CK(clk), .RN(n4238), .QN(n637) );
  DFFRX1 \block_r_reg[7][66]  ( .D(n2814), .CK(clk), .RN(n4238), .QN(n126) );
  DFFRX1 \block_r_reg[5][66]  ( .D(n3070), .CK(clk), .RN(n4238), .QN(n382) );
  DFFRX1 \block_r_reg[3][66]  ( .D(n3326), .CK(clk), .RN(n4238), .QN(n638) );
  DFFRX1 \block_r_reg[7][65]  ( .D(n2815), .CK(clk), .RN(n4237), .QN(n127) );
  DFFRX1 \block_r_reg[5][65]  ( .D(n3071), .CK(clk), .RN(n4237), .QN(n383) );
  DFFRX1 \block_r_reg[3][65]  ( .D(n3327), .CK(clk), .RN(n4237), .QN(n639) );
  DFFRX1 \block_r_reg[7][64]  ( .D(n2816), .CK(clk), .RN(n4237), .QN(n128) );
  DFFRX1 \block_r_reg[5][64]  ( .D(n3072), .CK(clk), .RN(n4237), .QN(n384) );
  DFFRX1 \block_r_reg[3][64]  ( .D(n3328), .CK(clk), .RN(n4236), .QN(n640) );
  DFFRX1 \block_r_reg[7][63]  ( .D(n2817), .CK(clk), .RN(n4236), .QN(n129) );
  DFFRX1 \block_r_reg[5][63]  ( .D(n3073), .CK(clk), .RN(n4236), .QN(n385) );
  DFFRX1 \block_r_reg[3][63]  ( .D(n3329), .CK(clk), .RN(n4236), .QN(n641) );
  DFFRX1 \block_r_reg[7][62]  ( .D(n2818), .CK(clk), .RN(n4235), .QN(n130) );
  DFFRX1 \block_r_reg[5][62]  ( .D(n3074), .CK(clk), .RN(n4235), .QN(n386) );
  DFFRX1 \block_r_reg[3][62]  ( .D(n3330), .CK(clk), .RN(n4235), .QN(n642) );
  DFFRX1 \block_r_reg[7][61]  ( .D(n2819), .CK(clk), .RN(n4235), .QN(n131) );
  DFFRX1 \block_r_reg[5][61]  ( .D(n3075), .CK(clk), .RN(n4235), .QN(n387) );
  DFFRX1 \block_r_reg[3][61]  ( .D(n3331), .CK(clk), .RN(n4234), .QN(n643) );
  DFFRX1 \block_r_reg[7][60]  ( .D(n2820), .CK(clk), .RN(n4234), .QN(n132) );
  DFFRX1 \block_r_reg[5][60]  ( .D(n3076), .CK(clk), .RN(n4234), .QN(n388) );
  DFFRX1 \block_r_reg[3][60]  ( .D(n3332), .CK(clk), .RN(n4234), .QN(n644) );
  DFFRX1 \block_r_reg[7][59]  ( .D(n2821), .CK(clk), .RN(n4233), .QN(n133) );
  DFFRX1 \block_r_reg[5][59]  ( .D(n3077), .CK(clk), .RN(n4233), .QN(n389) );
  DFFRX1 \block_r_reg[3][59]  ( .D(n3333), .CK(clk), .RN(n4233), .QN(n645) );
  DFFRX1 \block_r_reg[7][58]  ( .D(n2822), .CK(clk), .RN(n4233), .QN(n134) );
  DFFRX1 \block_r_reg[5][58]  ( .D(n3078), .CK(clk), .RN(n4233), .QN(n390) );
  DFFRX1 \block_r_reg[3][58]  ( .D(n3334), .CK(clk), .RN(n4232), .QN(n646) );
  DFFRX1 \block_r_reg[7][57]  ( .D(n2823), .CK(clk), .RN(n4232), .QN(n135) );
  DFFRX1 \block_r_reg[5][57]  ( .D(n3079), .CK(clk), .RN(n4232), .QN(n391) );
  DFFRX1 \block_r_reg[3][57]  ( .D(n3335), .CK(clk), .RN(n4232), .QN(n647) );
  DFFRX1 \block_r_reg[7][56]  ( .D(n2824), .CK(clk), .RN(n4231), .QN(n136) );
  DFFRX1 \block_r_reg[5][56]  ( .D(n3080), .CK(clk), .RN(n4231), .QN(n392) );
  DFFRX1 \block_r_reg[3][56]  ( .D(n3336), .CK(clk), .RN(n4231), .QN(n648) );
  DFFRX1 \block_r_reg[7][55]  ( .D(n2825), .CK(clk), .RN(n4231), .QN(n137) );
  DFFRX1 \block_r_reg[5][55]  ( .D(n3081), .CK(clk), .RN(n4231), .QN(n393) );
  DFFRX1 \block_r_reg[3][55]  ( .D(n3337), .CK(clk), .RN(n4230), .QN(n649) );
  DFFRX1 \block_r_reg[7][54]  ( .D(n2826), .CK(clk), .RN(n4230), .QN(n138) );
  DFFRX1 \block_r_reg[5][54]  ( .D(n3082), .CK(clk), .RN(n4230), .QN(n394) );
  DFFRX1 \block_r_reg[3][54]  ( .D(n3338), .CK(clk), .RN(n4230), .QN(n650) );
  DFFRX1 \block_r_reg[7][53]  ( .D(n2827), .CK(clk), .RN(n4229), .QN(n139) );
  DFFRX1 \block_r_reg[5][53]  ( .D(n3083), .CK(clk), .RN(n4229), .QN(n395) );
  DFFRX1 \block_r_reg[3][53]  ( .D(n3339), .CK(clk), .RN(n4229), .QN(n651) );
  DFFRX1 \block_r_reg[7][52]  ( .D(n2828), .CK(clk), .RN(n4229), .QN(n140) );
  DFFRX1 \block_r_reg[5][52]  ( .D(n3084), .CK(clk), .RN(n4229), .QN(n396) );
  DFFRX1 \block_r_reg[3][52]  ( .D(n3340), .CK(clk), .RN(n4228), .QN(n652) );
  DFFRX1 \block_r_reg[7][51]  ( .D(n2829), .CK(clk), .RN(n4228), .QN(n141) );
  DFFRX1 \block_r_reg[5][51]  ( .D(n3085), .CK(clk), .RN(n4228), .QN(n397) );
  DFFRX1 \block_r_reg[3][51]  ( .D(n3341), .CK(clk), .RN(n4228), .QN(n653) );
  DFFRX1 \block_r_reg[7][50]  ( .D(n2830), .CK(clk), .RN(n4227), .QN(n142) );
  DFFRX1 \block_r_reg[5][50]  ( .D(n3086), .CK(clk), .RN(n4227), .QN(n398) );
  DFFRX1 \block_r_reg[3][50]  ( .D(n3342), .CK(clk), .RN(n4227), .QN(n654) );
  DFFRX1 \block_r_reg[7][49]  ( .D(n2831), .CK(clk), .RN(n4227), .QN(n143) );
  DFFRX1 \block_r_reg[5][49]  ( .D(n3087), .CK(clk), .RN(n4227), .QN(n399) );
  DFFRX1 \block_r_reg[3][49]  ( .D(n3343), .CK(clk), .RN(n4226), .QN(n655) );
  DFFRX1 \block_r_reg[7][48]  ( .D(n2832), .CK(clk), .RN(n4226), .QN(n144) );
  DFFRX1 \block_r_reg[5][48]  ( .D(n3088), .CK(clk), .RN(n4226), .QN(n400) );
  DFFRX1 \block_r_reg[3][48]  ( .D(n3344), .CK(clk), .RN(n4226), .QN(n656) );
  DFFRX1 \block_r_reg[7][47]  ( .D(n2833), .CK(clk), .RN(n4225), .QN(n145) );
  DFFRX1 \block_r_reg[5][47]  ( .D(n3089), .CK(clk), .RN(n4225), .QN(n401) );
  DFFRX1 \block_r_reg[3][47]  ( .D(n3345), .CK(clk), .RN(n4225), .QN(n657) );
  DFFRX1 \block_r_reg[7][46]  ( .D(n2834), .CK(clk), .RN(n4225), .QN(n146) );
  DFFRX1 \block_r_reg[5][46]  ( .D(n3090), .CK(clk), .RN(n4225), .QN(n402) );
  DFFRX1 \block_r_reg[3][46]  ( .D(n3346), .CK(clk), .RN(n4224), .QN(n658) );
  DFFRX1 \block_r_reg[7][45]  ( .D(n2835), .CK(clk), .RN(n4224), .QN(n147) );
  DFFRX1 \block_r_reg[5][45]  ( .D(n3091), .CK(clk), .RN(n4224), .QN(n403) );
  DFFRX1 \block_r_reg[3][45]  ( .D(n3347), .CK(clk), .RN(n4224), .QN(n659) );
  DFFRX1 \block_r_reg[7][44]  ( .D(n2836), .CK(clk), .RN(n4223), .QN(n148) );
  DFFRX1 \block_r_reg[5][44]  ( .D(n3092), .CK(clk), .RN(n4223), .QN(n404) );
  DFFRX1 \block_r_reg[3][44]  ( .D(n3348), .CK(clk), .RN(n4223), .QN(n660) );
  DFFRX1 \block_r_reg[7][43]  ( .D(n2837), .CK(clk), .RN(n4223), .QN(n149) );
  DFFRX1 \block_r_reg[5][43]  ( .D(n3093), .CK(clk), .RN(n4223), .QN(n405) );
  DFFRX1 \block_r_reg[3][43]  ( .D(n3349), .CK(clk), .RN(n4222), .QN(n661) );
  DFFRX1 \block_r_reg[7][42]  ( .D(n2838), .CK(clk), .RN(n4222), .QN(n150) );
  DFFRX1 \block_r_reg[5][42]  ( .D(n3094), .CK(clk), .RN(n4222), .QN(n406) );
  DFFRX1 \block_r_reg[3][42]  ( .D(n3350), .CK(clk), .RN(n4222), .QN(n662) );
  DFFRX1 \block_r_reg[7][41]  ( .D(n2839), .CK(clk), .RN(n4221), .QN(n151) );
  DFFRX1 \block_r_reg[5][41]  ( .D(n3095), .CK(clk), .RN(n4221), .QN(n407) );
  DFFRX1 \block_r_reg[3][41]  ( .D(n3351), .CK(clk), .RN(n4221), .QN(n663) );
  DFFRX1 \block_r_reg[7][40]  ( .D(n2840), .CK(clk), .RN(n4221), .QN(n152) );
  DFFRX1 \block_r_reg[5][40]  ( .D(n3096), .CK(clk), .RN(n4221), .QN(n408) );
  DFFRX1 \block_r_reg[3][40]  ( .D(n3352), .CK(clk), .RN(n4220), .QN(n664) );
  DFFRX1 \block_r_reg[7][39]  ( .D(n2841), .CK(clk), .RN(n4220), .QN(n153) );
  DFFRX1 \block_r_reg[5][39]  ( .D(n3097), .CK(clk), .RN(n4220), .QN(n409) );
  DFFRX1 \block_r_reg[3][39]  ( .D(n3353), .CK(clk), .RN(n4220), .QN(n665) );
  DFFRX1 \block_r_reg[7][38]  ( .D(n2842), .CK(clk), .RN(n4219), .QN(n154) );
  DFFRX1 \block_r_reg[5][38]  ( .D(n3098), .CK(clk), .RN(n4219), .QN(n410) );
  DFFRX1 \block_r_reg[3][38]  ( .D(n3354), .CK(clk), .RN(n4219), .QN(n666) );
  DFFRX1 \block_r_reg[7][37]  ( .D(n2843), .CK(clk), .RN(n4219), .QN(n155) );
  DFFRX1 \block_r_reg[5][37]  ( .D(n3099), .CK(clk), .RN(n4219), .QN(n411) );
  DFFRX1 \block_r_reg[3][37]  ( .D(n3355), .CK(clk), .RN(n4218), .QN(n667) );
  DFFRX1 \block_r_reg[7][36]  ( .D(n2844), .CK(clk), .RN(n4218), .QN(n156) );
  DFFRX1 \block_r_reg[5][36]  ( .D(n3100), .CK(clk), .RN(n4218), .QN(n412) );
  DFFRX1 \block_r_reg[3][36]  ( .D(n3356), .CK(clk), .RN(n4218), .QN(n668) );
  DFFRX1 \block_r_reg[7][35]  ( .D(n2845), .CK(clk), .RN(n4217), .QN(n157) );
  DFFRX1 \block_r_reg[5][35]  ( .D(n3101), .CK(clk), .RN(n4217), .QN(n413) );
  DFFRX1 \block_r_reg[3][35]  ( .D(n3357), .CK(clk), .RN(n4217), .QN(n669) );
  DFFRX1 \block_r_reg[7][34]  ( .D(n2846), .CK(clk), .RN(n4217), .QN(n158) );
  DFFRX1 \block_r_reg[5][34]  ( .D(n3102), .CK(clk), .RN(n4217), .QN(n414) );
  DFFRX1 \block_r_reg[4][34]  ( .D(n3230), .CK(clk), .RN(n4216), .QN(n542) );
  DFFRX1 \block_r_reg[3][34]  ( .D(n3358), .CK(clk), .RN(n4216), .QN(n670) );
  DFFRX1 \block_r_reg[7][33]  ( .D(n2847), .CK(clk), .RN(n4216), .QN(n159) );
  DFFRX1 \block_r_reg[5][33]  ( .D(n3103), .CK(clk), .RN(n4216), .QN(n415) );
  DFFRX1 \block_r_reg[4][33]  ( .D(n3231), .CK(clk), .RN(n4216), .QN(n543) );
  DFFRX1 \block_r_reg[3][33]  ( .D(n3359), .CK(clk), .RN(n4216), .QN(n671) );
  DFFRX1 \block_r_reg[7][32]  ( .D(n2848), .CK(clk), .RN(n4215), .QN(n160) );
  DFFRX1 \block_r_reg[5][32]  ( .D(n3104), .CK(clk), .RN(n4215), .QN(n416) );
  DFFRX1 \block_r_reg[4][32]  ( .D(n3232), .CK(clk), .RN(n4215), .QN(n544) );
  DFFRX1 \block_r_reg[3][32]  ( .D(n3360), .CK(clk), .RN(n4215), .QN(n672) );
  DFFRX1 \block_r_reg[7][31]  ( .D(n2849), .CK(clk), .RN(n4215), .QN(n161) );
  DFFRX1 \block_r_reg[5][31]  ( .D(n3105), .CK(clk), .RN(n4215), .QN(n417) );
  DFFRX1 \block_r_reg[4][31]  ( .D(n3233), .CK(clk), .RN(n4214), .QN(n545) );
  DFFRX1 \block_r_reg[3][31]  ( .D(n3361), .CK(clk), .RN(n4214), .QN(n673) );
  DFFRX1 \block_r_reg[7][30]  ( .D(n2850), .CK(clk), .RN(n4214), .QN(n162) );
  DFFRX1 \block_r_reg[5][30]  ( .D(n3106), .CK(clk), .RN(n4214), .QN(n418) );
  DFFRX1 \block_r_reg[4][30]  ( .D(n3234), .CK(clk), .RN(n4214), .QN(n546) );
  DFFRX1 \block_r_reg[3][30]  ( .D(n3362), .CK(clk), .RN(n4214), .QN(n674) );
  DFFRX1 \block_r_reg[7][29]  ( .D(n2851), .CK(clk), .RN(n4213), .QN(n163) );
  DFFRX1 \block_r_reg[5][29]  ( .D(n3107), .CK(clk), .RN(n4213), .QN(n419) );
  DFFRX1 \block_r_reg[3][29]  ( .D(n3363), .CK(clk), .RN(n4213), .QN(n675) );
  DFFRX1 \block_r_reg[7][28]  ( .D(n2852), .CK(clk), .RN(n4213), .QN(n164) );
  DFFRX1 \block_r_reg[5][28]  ( .D(n3108), .CK(clk), .RN(n4213), .QN(n420) );
  DFFRX1 \block_r_reg[3][28]  ( .D(n3364), .CK(clk), .RN(n4212), .QN(n676) );
  DFFRX1 \block_r_reg[7][27]  ( .D(n2853), .CK(clk), .RN(n4212), .QN(n165) );
  DFFRX1 \block_r_reg[5][27]  ( .D(n3109), .CK(clk), .RN(n4212), .QN(n421) );
  DFFRX1 \block_r_reg[3][27]  ( .D(n3365), .CK(clk), .RN(n4212), .QN(n677) );
  DFFRX1 \block_r_reg[7][26]  ( .D(n2854), .CK(clk), .RN(n4211), .QN(n166) );
  DFFRX1 \block_r_reg[5][26]  ( .D(n3110), .CK(clk), .RN(n4211), .QN(n422) );
  DFFRX1 \block_r_reg[3][26]  ( .D(n3366), .CK(clk), .RN(n4211), .QN(n678) );
  DFFRX1 \block_r_reg[7][25]  ( .D(n2855), .CK(clk), .RN(n4211), .QN(n167) );
  DFFRX1 \block_r_reg[5][25]  ( .D(n3111), .CK(clk), .RN(n4211), .QN(n423) );
  DFFRX1 \block_r_reg[3][25]  ( .D(n3367), .CK(clk), .RN(n4210), .QN(n679) );
  DFFRX1 \block_r_reg[7][24]  ( .D(n2856), .CK(clk), .RN(n4210), .QN(n168) );
  DFFRX1 \block_r_reg[5][24]  ( .D(n3112), .CK(clk), .RN(n4210), .QN(n424) );
  DFFRX1 \block_r_reg[3][24]  ( .D(n3368), .CK(clk), .RN(n4210), .QN(n680) );
  DFFRX1 \block_r_reg[7][23]  ( .D(n2857), .CK(clk), .RN(n4209), .QN(n169) );
  DFFRX1 \block_r_reg[5][23]  ( .D(n3113), .CK(clk), .RN(n4209), .QN(n425) );
  DFFRX1 \block_r_reg[3][23]  ( .D(n3369), .CK(clk), .RN(n4209), .QN(n681) );
  DFFRX1 \block_r_reg[7][22]  ( .D(n2858), .CK(clk), .RN(n4209), .QN(n170) );
  DFFRX1 \block_r_reg[5][22]  ( .D(n3114), .CK(clk), .RN(n4209), .QN(n426) );
  DFFRX1 \block_r_reg[3][22]  ( .D(n3370), .CK(clk), .RN(n4208), .QN(n682) );
  DFFRX1 \block_r_reg[7][21]  ( .D(n2859), .CK(clk), .RN(n4208), .QN(n171) );
  DFFRX1 \block_r_reg[5][21]  ( .D(n3115), .CK(clk), .RN(n4208), .QN(n427) );
  DFFRX1 \block_r_reg[4][21]  ( .D(n3243), .CK(clk), .RN(n4208), .QN(n555) );
  DFFRX1 \block_r_reg[3][21]  ( .D(n3371), .CK(clk), .RN(n4208), .QN(n683) );
  DFFRX1 \block_r_reg[7][20]  ( .D(n2860), .CK(clk), .RN(n4207), .QN(n172) );
  DFFRX1 \block_r_reg[5][20]  ( .D(n3116), .CK(clk), .RN(n4207), .QN(n428) );
  DFFRX1 \block_r_reg[4][20]  ( .D(n3244), .CK(clk), .RN(n4207), .QN(n556) );
  DFFRX1 \block_r_reg[3][20]  ( .D(n3372), .CK(clk), .RN(n4207), .QN(n684) );
  DFFRX1 \block_r_reg[7][19]  ( .D(n2861), .CK(clk), .RN(n4207), .QN(n173) );
  DFFRX1 \block_r_reg[5][19]  ( .D(n3117), .CK(clk), .RN(n4207), .QN(n429) );
  DFFRX1 \block_r_reg[4][19]  ( .D(n3245), .CK(clk), .RN(n4206), .QN(n557) );
  DFFRX1 \block_r_reg[3][19]  ( .D(n3373), .CK(clk), .RN(n4206), .QN(n685) );
  DFFRX1 \block_r_reg[7][18]  ( .D(n2862), .CK(clk), .RN(n4206), .QN(n174) );
  DFFRX1 \block_r_reg[5][18]  ( .D(n3118), .CK(clk), .RN(n4206), .QN(n430) );
  DFFRX1 \block_r_reg[3][18]  ( .D(n3374), .CK(clk), .RN(n4206), .QN(n686) );
  DFFRX1 \block_r_reg[0][17]  ( .D(n3759), .CK(clk), .RN(n4291), .QN(n1071) );
  DFFRX1 \block_r_reg[6][17]  ( .D(n2991), .CK(clk), .RN(n4291), .QN(n303) );
  DFFRX1 \block_r_reg[4][17]  ( .D(n3247), .CK(clk), .RN(n4290), .QN(n559) );
  DFFRX1 \block_r_reg[2][17]  ( .D(n3503), .CK(clk), .RN(n4290), .QN(n815) );
  DFFRX1 \block_r_reg[0][16]  ( .D(n3760), .CK(clk), .RN(n4290), .QN(n1072) );
  DFFRX1 \block_r_reg[6][16]  ( .D(n2992), .CK(clk), .RN(n4290), .QN(n304) );
  DFFRX1 \block_r_reg[4][16]  ( .D(n3248), .CK(clk), .RN(n4290), .QN(n560) );
  DFFRX1 \block_r_reg[2][16]  ( .D(n3504), .CK(clk), .RN(n4290), .QN(n816) );
  DFFRX1 \block_r_reg[0][15]  ( .D(n3761), .CK(clk), .RN(n4289), .QN(n1073) );
  DFFRX1 \block_r_reg[6][15]  ( .D(n2993), .CK(clk), .RN(n4289), .QN(n305) );
  DFFRX1 \block_r_reg[4][15]  ( .D(n3249), .CK(clk), .RN(n4289), .QN(n561) );
  DFFRX1 \block_r_reg[2][15]  ( .D(n3505), .CK(clk), .RN(n4289), .QN(n817) );
  DFFRX1 \block_r_reg[0][14]  ( .D(n3762), .CK(clk), .RN(n4289), .QN(n1074) );
  DFFRX1 \block_r_reg[6][14]  ( .D(n2994), .CK(clk), .RN(n4289), .QN(n306) );
  DFFRX1 \block_r_reg[4][14]  ( .D(n3250), .CK(clk), .RN(n4288), .QN(n562) );
  DFFRX1 \block_r_reg[2][14]  ( .D(n3506), .CK(clk), .RN(n4288), .QN(n818) );
  DFFRX1 \block_r_reg[0][13]  ( .D(n3763), .CK(clk), .RN(n4288), .QN(n1075) );
  DFFRX1 \block_r_reg[6][13]  ( .D(n2995), .CK(clk), .RN(n4288), .QN(n307) );
  DFFRX1 \block_r_reg[4][13]  ( .D(n3251), .CK(clk), .RN(n4288), .QN(n563) );
  DFFRX1 \block_r_reg[2][13]  ( .D(n3507), .CK(clk), .RN(n4288), .QN(n819) );
  DFFRX1 \block_r_reg[0][12]  ( .D(n3764), .CK(clk), .RN(n4287), .QN(n1076) );
  DFFRX1 \block_r_reg[6][12]  ( .D(n2996), .CK(clk), .RN(n4287), .QN(n308) );
  DFFRX1 \block_r_reg[4][12]  ( .D(n3252), .CK(clk), .RN(n4287), .QN(n564) );
  DFFRX1 \block_r_reg[2][12]  ( .D(n3508), .CK(clk), .RN(n4287), .QN(n820) );
  DFFRX1 \block_r_reg[0][11]  ( .D(n3765), .CK(clk), .RN(n4287), .QN(n1077) );
  DFFRX1 \block_r_reg[6][11]  ( .D(n2997), .CK(clk), .RN(n4287), .QN(n309) );
  DFFRX1 \block_r_reg[4][11]  ( .D(n3253), .CK(clk), .RN(n4286), .QN(n565) );
  DFFRX1 \block_r_reg[2][11]  ( .D(n3509), .CK(clk), .RN(n4286), .QN(n821) );
  DFFRX1 \block_r_reg[0][10]  ( .D(n3766), .CK(clk), .RN(n4286), .QN(n1078) );
  DFFRX1 \block_r_reg[6][10]  ( .D(n2998), .CK(clk), .RN(n4286), .QN(n310) );
  DFFRX1 \block_r_reg[4][10]  ( .D(n3254), .CK(clk), .RN(n4286), .QN(n566) );
  DFFRX1 \block_r_reg[2][10]  ( .D(n3510), .CK(clk), .RN(n4286), .QN(n822) );
  DFFRX1 \block_r_reg[0][9]  ( .D(n3767), .CK(clk), .RN(n4285), .QN(n1079) );
  DFFRX1 \block_r_reg[6][9]  ( .D(n2999), .CK(clk), .RN(n4285), .QN(n311) );
  DFFRX1 \block_r_reg[4][9]  ( .D(n3255), .CK(clk), .RN(n4285), .QN(n567) );
  DFFRX1 \block_r_reg[2][9]  ( .D(n3511), .CK(clk), .RN(n4285), .QN(n823) );
  DFFRX1 \block_r_reg[0][8]  ( .D(n3768), .CK(clk), .RN(n4285), .QN(n1080) );
  DFFRX1 \block_r_reg[6][8]  ( .D(n3000), .CK(clk), .RN(n4285), .QN(n312) );
  DFFRX1 \block_r_reg[4][8]  ( .D(n3256), .CK(clk), .RN(n4284), .QN(n568) );
  DFFRX1 \block_r_reg[2][8]  ( .D(n3512), .CK(clk), .RN(n4284), .QN(n824) );
  DFFRX1 \block_r_reg[0][7]  ( .D(n3769), .CK(clk), .RN(n4284), .QN(n1081) );
  DFFRX1 \block_r_reg[6][7]  ( .D(n3001), .CK(clk), .RN(n4284), .QN(n313) );
  DFFRX1 \block_r_reg[4][7]  ( .D(n3257), .CK(clk), .RN(n4284), .QN(n569) );
  DFFRX1 \block_r_reg[2][7]  ( .D(n3513), .CK(clk), .RN(n4284), .QN(n825) );
  DFFRX1 \block_r_reg[0][6]  ( .D(n3770), .CK(clk), .RN(n4283), .QN(n1082) );
  DFFRX1 \block_r_reg[6][6]  ( .D(n3002), .CK(clk), .RN(n4283), .QN(n314) );
  DFFRX1 \block_r_reg[4][6]  ( .D(n3258), .CK(clk), .RN(n4283), .QN(n570) );
  DFFRX1 \block_r_reg[2][6]  ( .D(n3514), .CK(clk), .RN(n4283), .QN(n826) );
  DFFRX1 \block_r_reg[0][5]  ( .D(n3771), .CK(clk), .RN(n4283), .QN(n1083) );
  DFFRX1 \block_r_reg[6][5]  ( .D(n3003), .CK(clk), .RN(n4283), .QN(n315) );
  DFFRX1 \block_r_reg[4][5]  ( .D(n3259), .CK(clk), .RN(n4282), .QN(n571) );
  DFFRX1 \block_r_reg[2][5]  ( .D(n3515), .CK(clk), .RN(n4282), .QN(n827) );
  DFFRX1 \block_r_reg[0][4]  ( .D(n3772), .CK(clk), .RN(n4282), .QN(n1084) );
  DFFRX1 \block_r_reg[6][4]  ( .D(n3004), .CK(clk), .RN(n4282), .QN(n316) );
  DFFRX1 \block_r_reg[4][4]  ( .D(n3260), .CK(clk), .RN(n4282), .QN(n572) );
  DFFRX1 \block_r_reg[2][4]  ( .D(n3516), .CK(clk), .RN(n4282), .QN(n828) );
  DFFRX1 \block_r_reg[0][3]  ( .D(n3773), .CK(clk), .RN(n4281), .QN(n1085) );
  DFFRX1 \block_r_reg[6][3]  ( .D(n3005), .CK(clk), .RN(n4281), .QN(n317) );
  DFFRX1 \block_r_reg[4][3]  ( .D(n3261), .CK(clk), .RN(n4281), .QN(n573) );
  DFFRX1 \block_r_reg[2][3]  ( .D(n3517), .CK(clk), .RN(n4281), .QN(n829) );
  DFFRX1 \block_r_reg[0][2]  ( .D(n3774), .CK(clk), .RN(n4281), .QN(n1086) );
  DFFRX1 \block_r_reg[6][2]  ( .D(n3006), .CK(clk), .RN(n4281), .QN(n318) );
  DFFRX1 \block_r_reg[4][2]  ( .D(n3262), .CK(clk), .RN(n4280), .QN(n574) );
  DFFRX1 \block_r_reg[2][2]  ( .D(n3518), .CK(clk), .RN(n4280), .QN(n830) );
  DFFRX1 \block_r_reg[0][1]  ( .D(n3775), .CK(clk), .RN(n4280), .QN(n1087) );
  DFFRX1 \block_r_reg[6][1]  ( .D(n3007), .CK(clk), .RN(n4280), .QN(n319) );
  DFFRX1 \block_r_reg[4][1]  ( .D(n3263), .CK(clk), .RN(n4280), .QN(n575) );
  DFFRX1 \block_r_reg[2][1]  ( .D(n3519), .CK(clk), .RN(n4280), .QN(n831) );
  DFFRX1 \block_r_reg[0][0]  ( .D(n3776), .CK(clk), .RN(n4279), .QN(n1088) );
  DFFRX1 \block_r_reg[6][0]  ( .D(n3008), .CK(clk), .RN(n4279), .QN(n320) );
  DFFRX1 \block_r_reg[4][0]  ( .D(n3264), .CK(clk), .RN(n4279), .QN(n576) );
  DFFRX1 \block_r_reg[2][0]  ( .D(n3520), .CK(clk), .RN(n4279), .QN(n832) );
  DFFRX1 \block_r_reg[0][127]  ( .D(n3649), .CK(clk), .RN(n4279), .QN(n961) );
  DFFRX1 \block_r_reg[6][127]  ( .D(n2881), .CK(clk), .RN(n4279), .QN(n193) );
  DFFRX1 \block_r_reg[2][127]  ( .D(n3393), .CK(clk), .RN(n4278), .QN(n705) );
  DFFRX1 \block_r_reg[0][126]  ( .D(n3650), .CK(clk), .RN(n4278), .QN(n962) );
  DFFRX1 \block_r_reg[6][126]  ( .D(n2882), .CK(clk), .RN(n4278), .QN(n194) );
  DFFRX1 \block_r_reg[2][126]  ( .D(n3394), .CK(clk), .RN(n4278), .QN(n706) );
  DFFRX1 \block_r_reg[0][125]  ( .D(n3651), .CK(clk), .RN(n4277), .QN(n963) );
  DFFRX1 \block_r_reg[6][125]  ( .D(n2883), .CK(clk), .RN(n4277), .QN(n195) );
  DFFRX1 \block_r_reg[2][125]  ( .D(n3395), .CK(clk), .RN(n4277), .QN(n707) );
  DFFRX1 \block_r_reg[0][124]  ( .D(n3652), .CK(clk), .RN(n4277), .QN(n964) );
  DFFRX1 \block_r_reg[6][124]  ( .D(n2884), .CK(clk), .RN(n4277), .QN(n196) );
  DFFRX1 \block_r_reg[2][124]  ( .D(n3396), .CK(clk), .RN(n4276), .QN(n708) );
  DFFRX1 \block_r_reg[0][123]  ( .D(n3653), .CK(clk), .RN(n4276), .QN(n965) );
  DFFRX1 \block_r_reg[6][123]  ( .D(n2885), .CK(clk), .RN(n4276), .QN(n197) );
  DFFRX1 \block_r_reg[2][123]  ( .D(n3397), .CK(clk), .RN(n4276), .QN(n709) );
  DFFRX1 \block_r_reg[0][122]  ( .D(n3654), .CK(clk), .RN(n4275), .QN(n966) );
  DFFRX1 \block_r_reg[6][122]  ( .D(n2886), .CK(clk), .RN(n4275), .QN(n198) );
  DFFRX1 \block_r_reg[2][122]  ( .D(n3398), .CK(clk), .RN(n4275), .QN(n710) );
  DFFRX1 \block_r_reg[0][121]  ( .D(n3655), .CK(clk), .RN(n4275), .QN(n967) );
  DFFRX1 \block_r_reg[6][121]  ( .D(n2887), .CK(clk), .RN(n4275), .QN(n199) );
  DFFRX1 \block_r_reg[2][121]  ( .D(n3399), .CK(clk), .RN(n4274), .QN(n711) );
  DFFRX1 \block_r_reg[0][120]  ( .D(n3656), .CK(clk), .RN(n4274), .QN(n968) );
  DFFRX1 \block_r_reg[6][120]  ( .D(n2888), .CK(clk), .RN(n4274), .QN(n200) );
  DFFRX1 \block_r_reg[2][120]  ( .D(n3400), .CK(clk), .RN(n4274), .QN(n712) );
  DFFRX1 \block_r_reg[0][119]  ( .D(n3657), .CK(clk), .RN(n4273), .QN(n969) );
  DFFRX1 \block_r_reg[6][119]  ( .D(n2889), .CK(clk), .RN(n4273), .QN(n201) );
  DFFRX1 \block_r_reg[2][119]  ( .D(n3401), .CK(clk), .RN(n4273), .QN(n713) );
  DFFRX1 \block_r_reg[0][118]  ( .D(n3658), .CK(clk), .RN(n4273), .QN(n970) );
  DFFRX1 \block_r_reg[6][118]  ( .D(n2890), .CK(clk), .RN(n4273), .QN(n202) );
  DFFRX1 \block_r_reg[2][118]  ( .D(n3402), .CK(clk), .RN(n4272), .QN(n714) );
  DFFRX1 \block_r_reg[0][117]  ( .D(n3659), .CK(clk), .RN(n4272), .QN(n971) );
  DFFRX1 \block_r_reg[6][117]  ( .D(n2891), .CK(clk), .RN(n4272), .QN(n203) );
  DFFRX1 \block_r_reg[4][117]  ( .D(n3147), .CK(clk), .RN(n4272), .QN(n459) );
  DFFRX1 \block_r_reg[2][117]  ( .D(n3403), .CK(clk), .RN(n4272), .QN(n715) );
  DFFRX1 \block_r_reg[0][116]  ( .D(n3660), .CK(clk), .RN(n4271), .QN(n972) );
  DFFRX1 \block_r_reg[6][116]  ( .D(n2892), .CK(clk), .RN(n4271), .QN(n204) );
  DFFRX1 \block_r_reg[4][116]  ( .D(n3148), .CK(clk), .RN(n4271), .QN(n460) );
  DFFRX1 \block_r_reg[2][116]  ( .D(n3404), .CK(clk), .RN(n4271), .QN(n716) );
  DFFRX1 \block_r_reg[0][115]  ( .D(n3661), .CK(clk), .RN(n4271), .QN(n973) );
  DFFRX1 \block_r_reg[6][115]  ( .D(n2893), .CK(clk), .RN(n4271), .QN(n205) );
  DFFRX1 \block_r_reg[4][115]  ( .D(n3149), .CK(clk), .RN(n4270), .QN(n461) );
  DFFRX1 \block_r_reg[2][115]  ( .D(n3405), .CK(clk), .RN(n4270), .QN(n717) );
  DFFRX1 \block_r_reg[0][114]  ( .D(n3662), .CK(clk), .RN(n4270), .QN(n974) );
  DFFRX1 \block_r_reg[6][114]  ( .D(n2894), .CK(clk), .RN(n4270), .QN(n206) );
  DFFRX1 \block_r_reg[4][114]  ( .D(n3150), .CK(clk), .RN(n4270), .QN(n462) );
  DFFRX1 \block_r_reg[2][114]  ( .D(n3406), .CK(clk), .RN(n4270), .QN(n718) );
  DFFRX1 \block_r_reg[0][113]  ( .D(n3663), .CK(clk), .RN(n4269), .QN(n975) );
  DFFRX1 \block_r_reg[6][113]  ( .D(n2895), .CK(clk), .RN(n4269), .QN(n207) );
  DFFRX1 \block_r_reg[4][113]  ( .D(n3151), .CK(clk), .RN(n4269), .QN(n463) );
  DFFRX1 \block_r_reg[2][113]  ( .D(n3407), .CK(clk), .RN(n4269), .QN(n719) );
  DFFRX1 \block_r_reg[0][112]  ( .D(n3664), .CK(clk), .RN(n4269), .QN(n976) );
  DFFRX1 \block_r_reg[6][112]  ( .D(n2896), .CK(clk), .RN(n4269), .QN(n208) );
  DFFRX1 \block_r_reg[4][112]  ( .D(n3152), .CK(clk), .RN(n4268), .QN(n464) );
  DFFRX1 \block_r_reg[2][112]  ( .D(n3408), .CK(clk), .RN(n4268), .QN(n720) );
  DFFRX1 \block_r_reg[0][111]  ( .D(n3665), .CK(clk), .RN(n4268), .QN(n977) );
  DFFRX1 \block_r_reg[6][111]  ( .D(n2897), .CK(clk), .RN(n4268), .QN(n209) );
  DFFRX1 \block_r_reg[4][111]  ( .D(n3153), .CK(clk), .RN(n4268), .QN(n465) );
  DFFRX1 \block_r_reg[2][111]  ( .D(n3409), .CK(clk), .RN(n4268), .QN(n721) );
  DFFRX1 \block_r_reg[0][110]  ( .D(n3666), .CK(clk), .RN(n4267), .QN(n978) );
  DFFRX1 \block_r_reg[6][110]  ( .D(n2898), .CK(clk), .RN(n4267), .QN(n210) );
  DFFRX1 \block_r_reg[4][110]  ( .D(n3154), .CK(clk), .RN(n4267), .QN(n466) );
  DFFRX1 \block_r_reg[2][110]  ( .D(n3410), .CK(clk), .RN(n4267), .QN(n722) );
  DFFRX1 \block_r_reg[0][109]  ( .D(n3667), .CK(clk), .RN(n4267), .QN(n979) );
  DFFRX1 \block_r_reg[6][109]  ( .D(n2899), .CK(clk), .RN(n4267), .QN(n211) );
  DFFRX1 \block_r_reg[4][109]  ( .D(n3155), .CK(clk), .RN(n4266), .QN(n467) );
  DFFRX1 \block_r_reg[2][109]  ( .D(n3411), .CK(clk), .RN(n4266), .QN(n723) );
  DFFRX1 \block_r_reg[0][108]  ( .D(n3668), .CK(clk), .RN(n4266), .QN(n980) );
  DFFRX1 \block_r_reg[6][108]  ( .D(n2900), .CK(clk), .RN(n4266), .QN(n212) );
  DFFRX1 \block_r_reg[4][108]  ( .D(n3156), .CK(clk), .RN(n4266), .QN(n468) );
  DFFRX1 \block_r_reg[2][108]  ( .D(n3412), .CK(clk), .RN(n4266), .QN(n724) );
  DFFRX1 \block_r_reg[0][107]  ( .D(n3669), .CK(clk), .RN(n4265), .QN(n981) );
  DFFRX1 \block_r_reg[6][107]  ( .D(n2901), .CK(clk), .RN(n4265), .QN(n213) );
  DFFRX1 \block_r_reg[4][107]  ( .D(n3157), .CK(clk), .RN(n4265), .QN(n469) );
  DFFRX1 \block_r_reg[2][107]  ( .D(n3413), .CK(clk), .RN(n4265), .QN(n725) );
  DFFRX1 \block_r_reg[0][106]  ( .D(n3670), .CK(clk), .RN(n4265), .QN(n982) );
  DFFRX1 \block_r_reg[6][106]  ( .D(n2902), .CK(clk), .RN(n4265), .QN(n214) );
  DFFRX1 \block_r_reg[4][106]  ( .D(n3158), .CK(clk), .RN(n4264), .QN(n470) );
  DFFRX1 \block_r_reg[2][106]  ( .D(n3414), .CK(clk), .RN(n4264), .QN(n726) );
  DFFRX1 \block_r_reg[0][105]  ( .D(n3671), .CK(clk), .RN(n4264), .QN(n983) );
  DFFRX1 \block_r_reg[6][105]  ( .D(n2903), .CK(clk), .RN(n4264), .QN(n215) );
  DFFRX1 \block_r_reg[4][105]  ( .D(n3159), .CK(clk), .RN(n4264), .QN(n471) );
  DFFRX1 \block_r_reg[2][105]  ( .D(n3415), .CK(clk), .RN(n4264), .QN(n727) );
  DFFRX1 \block_r_reg[0][104]  ( .D(n3672), .CK(clk), .RN(n4263), .QN(n984) );
  DFFRX1 \block_r_reg[6][104]  ( .D(n2904), .CK(clk), .RN(n4263), .QN(n216) );
  DFFRX1 \block_r_reg[4][104]  ( .D(n3160), .CK(clk), .RN(n4263), .QN(n472) );
  DFFRX1 \block_r_reg[2][104]  ( .D(n3416), .CK(clk), .RN(n4263), .QN(n728) );
  DFFRX1 \block_r_reg[0][103]  ( .D(n3673), .CK(clk), .RN(n4263), .QN(n985) );
  DFFRX1 \block_r_reg[6][103]  ( .D(n2905), .CK(clk), .RN(n4263), .QN(n217) );
  DFFRX1 \block_r_reg[4][103]  ( .D(n3161), .CK(clk), .RN(n4262), .QN(n473) );
  DFFRX1 \block_r_reg[2][103]  ( .D(n3417), .CK(clk), .RN(n4262), .QN(n729) );
  DFFRX1 \block_r_reg[0][102]  ( .D(n3674), .CK(clk), .RN(n4262), .QN(n986) );
  DFFRX1 \block_r_reg[6][102]  ( .D(n2906), .CK(clk), .RN(n4262), .QN(n218) );
  DFFRX1 \block_r_reg[4][102]  ( .D(n3162), .CK(clk), .RN(n4262), .QN(n474) );
  DFFRX1 \block_r_reg[2][102]  ( .D(n3418), .CK(clk), .RN(n4262), .QN(n730) );
  DFFRX1 \block_r_reg[0][101]  ( .D(n3675), .CK(clk), .RN(n4261), .QN(n987) );
  DFFRX1 \block_r_reg[6][101]  ( .D(n2907), .CK(clk), .RN(n4261), .QN(n219) );
  DFFRX1 \block_r_reg[4][101]  ( .D(n3163), .CK(clk), .RN(n4261), .QN(n475) );
  DFFRX1 \block_r_reg[2][101]  ( .D(n3419), .CK(clk), .RN(n4261), .QN(n731) );
  DFFRX1 \block_r_reg[0][100]  ( .D(n3676), .CK(clk), .RN(n4261), .QN(n988) );
  DFFRX1 \block_r_reg[6][100]  ( .D(n2908), .CK(clk), .RN(n4261), .QN(n220) );
  DFFRX1 \block_r_reg[4][100]  ( .D(n3164), .CK(clk), .RN(n4260), .QN(n476) );
  DFFRX1 \block_r_reg[2][100]  ( .D(n3420), .CK(clk), .RN(n4260), .QN(n732) );
  DFFRX1 \block_r_reg[0][99]  ( .D(n3677), .CK(clk), .RN(n4260), .QN(n989) );
  DFFRX1 \block_r_reg[6][99]  ( .D(n2909), .CK(clk), .RN(n4260), .QN(n221) );
  DFFRX1 \block_r_reg[4][99]  ( .D(n3165), .CK(clk), .RN(n4260), .QN(n477) );
  DFFRX1 \block_r_reg[2][99]  ( .D(n3421), .CK(clk), .RN(n4260), .QN(n733) );
  DFFRX1 \block_r_reg[0][98]  ( .D(n3678), .CK(clk), .RN(n4259), .QN(n990) );
  DFFRX1 \block_r_reg[6][98]  ( .D(n2910), .CK(clk), .RN(n4259), .QN(n222) );
  DFFRX1 \block_r_reg[4][98]  ( .D(n3166), .CK(clk), .RN(n4259), .QN(n478) );
  DFFRX1 \block_r_reg[2][98]  ( .D(n3422), .CK(clk), .RN(n4259), .QN(n734) );
  DFFRX1 \block_r_reg[0][97]  ( .D(n3679), .CK(clk), .RN(n4259), .QN(n991) );
  DFFRX1 \block_r_reg[6][97]  ( .D(n2911), .CK(clk), .RN(n4259), .QN(n223) );
  DFFRX1 \block_r_reg[4][97]  ( .D(n3167), .CK(clk), .RN(n4258), .QN(n479) );
  DFFRX1 \block_r_reg[2][97]  ( .D(n3423), .CK(clk), .RN(n4258), .QN(n735) );
  DFFRX1 \block_r_reg[0][96]  ( .D(n3680), .CK(clk), .RN(n4258), .QN(n992) );
  DFFRX1 \block_r_reg[6][96]  ( .D(n2912), .CK(clk), .RN(n4258), .QN(n224) );
  DFFRX1 \block_r_reg[4][96]  ( .D(n3168), .CK(clk), .RN(n4258), .QN(n480) );
  DFFRX1 \block_r_reg[2][96]  ( .D(n3424), .CK(clk), .RN(n4258), .QN(n736) );
  DFFRX1 \block_r_reg[0][95]  ( .D(n3681), .CK(clk), .RN(n4257), .QN(n993) );
  DFFRX1 \block_r_reg[6][95]  ( .D(n2913), .CK(clk), .RN(n4257), .QN(n225) );
  DFFRX1 \block_r_reg[4][95]  ( .D(n3169), .CK(clk), .RN(n4257), .QN(n481) );
  DFFRX1 \block_r_reg[2][95]  ( .D(n3425), .CK(clk), .RN(n4257), .QN(n737) );
  DFFRX1 \block_r_reg[0][94]  ( .D(n3682), .CK(clk), .RN(n4257), .QN(n994) );
  DFFRX1 \block_r_reg[6][94]  ( .D(n2914), .CK(clk), .RN(n4257), .QN(n226) );
  DFFRX1 \block_r_reg[4][94]  ( .D(n3170), .CK(clk), .RN(n4256), .QN(n482) );
  DFFRX1 \block_r_reg[2][94]  ( .D(n3426), .CK(clk), .RN(n4256), .QN(n738) );
  DFFRX1 \block_r_reg[0][93]  ( .D(n3683), .CK(clk), .RN(n4256), .QN(n995) );
  DFFRX1 \block_r_reg[6][93]  ( .D(n2915), .CK(clk), .RN(n4256), .QN(n227) );
  DFFRX1 \block_r_reg[4][93]  ( .D(n3171), .CK(clk), .RN(n4256), .QN(n483) );
  DFFRX1 \block_r_reg[2][93]  ( .D(n3427), .CK(clk), .RN(n4256), .QN(n739) );
  DFFRX1 \block_r_reg[0][92]  ( .D(n3684), .CK(clk), .RN(n4255), .QN(n996) );
  DFFRX1 \block_r_reg[6][92]  ( .D(n2916), .CK(clk), .RN(n4255), .QN(n228) );
  DFFRX1 \block_r_reg[4][92]  ( .D(n3172), .CK(clk), .RN(n4255), .QN(n484) );
  DFFRX1 \block_r_reg[2][92]  ( .D(n3428), .CK(clk), .RN(n4255), .QN(n740) );
  DFFRX1 \block_r_reg[0][91]  ( .D(n3685), .CK(clk), .RN(n4255), .QN(n997) );
  DFFRX1 \block_r_reg[6][91]  ( .D(n2917), .CK(clk), .RN(n4255), .QN(n229) );
  DFFRX1 \block_r_reg[4][91]  ( .D(n3173), .CK(clk), .RN(n4254), .QN(n485) );
  DFFRX1 \block_r_reg[2][91]  ( .D(n3429), .CK(clk), .RN(n4254), .QN(n741) );
  DFFRX1 \block_r_reg[0][90]  ( .D(n3686), .CK(clk), .RN(n4254), .QN(n998) );
  DFFRX1 \block_r_reg[6][90]  ( .D(n2918), .CK(clk), .RN(n4254), .QN(n230) );
  DFFRX1 \block_r_reg[4][90]  ( .D(n3174), .CK(clk), .RN(n4254), .QN(n486) );
  DFFRX1 \block_r_reg[2][90]  ( .D(n3430), .CK(clk), .RN(n4254), .QN(n742) );
  DFFRX1 \block_r_reg[0][89]  ( .D(n3687), .CK(clk), .RN(n4253), .QN(n999) );
  DFFRX1 \block_r_reg[6][89]  ( .D(n2919), .CK(clk), .RN(n4253), .QN(n231) );
  DFFRX1 \block_r_reg[4][89]  ( .D(n3175), .CK(clk), .RN(n4253), .QN(n487) );
  DFFRX1 \block_r_reg[2][89]  ( .D(n3431), .CK(clk), .RN(n4253), .QN(n743) );
  DFFRX1 \block_r_reg[0][88]  ( .D(n3688), .CK(clk), .RN(n4253), .QN(n1000) );
  DFFRX1 \block_r_reg[6][88]  ( .D(n2920), .CK(clk), .RN(n4253), .QN(n232) );
  DFFRX1 \block_r_reg[4][88]  ( .D(n3176), .CK(clk), .RN(n4252), .QN(n488) );
  DFFRX1 \block_r_reg[2][88]  ( .D(n3432), .CK(clk), .RN(n4252), .QN(n744) );
  DFFRX1 \block_r_reg[0][87]  ( .D(n3689), .CK(clk), .RN(n4252), .QN(n1001) );
  DFFRX1 \block_r_reg[6][87]  ( .D(n2921), .CK(clk), .RN(n4252), .QN(n233) );
  DFFRX1 \block_r_reg[4][87]  ( .D(n3177), .CK(clk), .RN(n4252), .QN(n489) );
  DFFRX1 \block_r_reg[2][87]  ( .D(n3433), .CK(clk), .RN(n4252), .QN(n745) );
  DFFRX1 \block_r_reg[0][86]  ( .D(n3690), .CK(clk), .RN(n4251), .QN(n1002) );
  DFFRX1 \block_r_reg[6][86]  ( .D(n2922), .CK(clk), .RN(n4251), .QN(n234) );
  DFFRX1 \block_r_reg[4][86]  ( .D(n3178), .CK(clk), .RN(n4251), .QN(n490) );
  DFFRX1 \block_r_reg[2][86]  ( .D(n3434), .CK(clk), .RN(n4251), .QN(n746) );
  DFFRX1 \block_r_reg[0][85]  ( .D(n3691), .CK(clk), .RN(n4251), .QN(n1003) );
  DFFRX1 \block_r_reg[6][85]  ( .D(n2923), .CK(clk), .RN(n4251), .QN(n235) );
  DFFRX1 \block_r_reg[4][85]  ( .D(n3179), .CK(clk), .RN(n4250), .QN(n491) );
  DFFRX1 \block_r_reg[2][85]  ( .D(n3435), .CK(clk), .RN(n4250), .QN(n747) );
  DFFRX1 \block_r_reg[0][84]  ( .D(n3692), .CK(clk), .RN(n4250), .QN(n1004) );
  DFFRX1 \block_r_reg[6][84]  ( .D(n2924), .CK(clk), .RN(n4250), .QN(n236) );
  DFFRX1 \block_r_reg[4][84]  ( .D(n3180), .CK(clk), .RN(n4250), .QN(n492) );
  DFFRX1 \block_r_reg[2][84]  ( .D(n3436), .CK(clk), .RN(n4250), .QN(n748) );
  DFFRX1 \block_r_reg[0][83]  ( .D(n3693), .CK(clk), .RN(n4249), .QN(n1005) );
  DFFRX1 \block_r_reg[6][83]  ( .D(n2925), .CK(clk), .RN(n4249), .QN(n237) );
  DFFRX1 \block_r_reg[4][83]  ( .D(n3181), .CK(clk), .RN(n4249), .QN(n493) );
  DFFRX1 \block_r_reg[2][83]  ( .D(n3437), .CK(clk), .RN(n4249), .QN(n749) );
  DFFRX1 \block_r_reg[0][82]  ( .D(n3694), .CK(clk), .RN(n4249), .QN(n1006) );
  DFFRX1 \block_r_reg[6][82]  ( .D(n2926), .CK(clk), .RN(n4249), .QN(n238) );
  DFFRX1 \block_r_reg[4][82]  ( .D(n3182), .CK(clk), .RN(n4248), .QN(n494) );
  DFFRX1 \block_r_reg[2][82]  ( .D(n3438), .CK(clk), .RN(n4248), .QN(n750) );
  DFFRX1 \block_r_reg[0][81]  ( .D(n3695), .CK(clk), .RN(n4248), .QN(n1007) );
  DFFRX1 \block_r_reg[6][81]  ( .D(n2927), .CK(clk), .RN(n4248), .QN(n239) );
  DFFRX1 \block_r_reg[4][81]  ( .D(n3183), .CK(clk), .RN(n4248), .QN(n495) );
  DFFRX1 \block_r_reg[2][81]  ( .D(n3439), .CK(clk), .RN(n4248), .QN(n751) );
  DFFRX1 \block_r_reg[0][80]  ( .D(n3696), .CK(clk), .RN(n4247), .QN(n1008) );
  DFFRX1 \block_r_reg[6][80]  ( .D(n2928), .CK(clk), .RN(n4247), .QN(n240) );
  DFFRX1 \block_r_reg[4][80]  ( .D(n3184), .CK(clk), .RN(n4247), .QN(n496) );
  DFFRX1 \block_r_reg[2][80]  ( .D(n3440), .CK(clk), .RN(n4247), .QN(n752) );
  DFFRX1 \block_r_reg[0][79]  ( .D(n3697), .CK(clk), .RN(n4247), .QN(n1009) );
  DFFRX1 \block_r_reg[6][79]  ( .D(n2929), .CK(clk), .RN(n4247), .QN(n241) );
  DFFRX1 \block_r_reg[4][79]  ( .D(n3185), .CK(clk), .RN(n4246), .QN(n497) );
  DFFRX1 \block_r_reg[2][79]  ( .D(n3441), .CK(clk), .RN(n4246), .QN(n753) );
  DFFRX1 \block_r_reg[0][78]  ( .D(n3698), .CK(clk), .RN(n4246), .QN(n1010) );
  DFFRX1 \block_r_reg[6][78]  ( .D(n2930), .CK(clk), .RN(n4246), .QN(n242) );
  DFFRX1 \block_r_reg[4][78]  ( .D(n3186), .CK(clk), .RN(n4246), .QN(n498) );
  DFFRX1 \block_r_reg[2][78]  ( .D(n3442), .CK(clk), .RN(n4246), .QN(n754) );
  DFFRX1 \block_r_reg[0][77]  ( .D(n3699), .CK(clk), .RN(n4245), .QN(n1011) );
  DFFRX1 \block_r_reg[6][77]  ( .D(n2931), .CK(clk), .RN(n4245), .QN(n243) );
  DFFRX1 \block_r_reg[4][77]  ( .D(n3187), .CK(clk), .RN(n4245), .QN(n499) );
  DFFRX1 \block_r_reg[2][77]  ( .D(n3443), .CK(clk), .RN(n4245), .QN(n755) );
  DFFRX1 \block_r_reg[0][76]  ( .D(n3700), .CK(clk), .RN(n4245), .QN(n1012) );
  DFFRX1 \block_r_reg[6][76]  ( .D(n2932), .CK(clk), .RN(n4245), .QN(n244) );
  DFFRX1 \block_r_reg[4][76]  ( .D(n3188), .CK(clk), .RN(n4244), .QN(n500) );
  DFFRX1 \block_r_reg[2][76]  ( .D(n3444), .CK(clk), .RN(n4244), .QN(n756) );
  DFFRX1 \block_r_reg[0][75]  ( .D(n3701), .CK(clk), .RN(n4244), .QN(n1013) );
  DFFRX1 \block_r_reg[6][75]  ( .D(n2933), .CK(clk), .RN(n4244), .QN(n245) );
  DFFRX1 \block_r_reg[4][75]  ( .D(n3189), .CK(clk), .RN(n4244), .QN(n501) );
  DFFRX1 \block_r_reg[2][75]  ( .D(n3445), .CK(clk), .RN(n4244), .QN(n757) );
  DFFRX1 \block_r_reg[0][74]  ( .D(n3702), .CK(clk), .RN(n4243), .QN(n1014) );
  DFFRX1 \block_r_reg[6][74]  ( .D(n2934), .CK(clk), .RN(n4243), .QN(n246) );
  DFFRX1 \block_r_reg[4][74]  ( .D(n3190), .CK(clk), .RN(n4243), .QN(n502) );
  DFFRX1 \block_r_reg[2][74]  ( .D(n3446), .CK(clk), .RN(n4243), .QN(n758) );
  DFFRX1 \block_r_reg[0][73]  ( .D(n3703), .CK(clk), .RN(n4243), .QN(n1015) );
  DFFRX1 \block_r_reg[6][73]  ( .D(n2935), .CK(clk), .RN(n4243), .QN(n247) );
  DFFRX1 \block_r_reg[4][73]  ( .D(n3191), .CK(clk), .RN(n4242), .QN(n503) );
  DFFRX1 \block_r_reg[2][73]  ( .D(n3447), .CK(clk), .RN(n4242), .QN(n759) );
  DFFRX1 \block_r_reg[0][72]  ( .D(n3704), .CK(clk), .RN(n4242), .QN(n1016) );
  DFFRX1 \block_r_reg[6][72]  ( .D(n2936), .CK(clk), .RN(n4242), .QN(n248) );
  DFFRX1 \block_r_reg[4][72]  ( .D(n3192), .CK(clk), .RN(n4242), .QN(n504) );
  DFFRX1 \block_r_reg[2][72]  ( .D(n3448), .CK(clk), .RN(n4242), .QN(n760) );
  DFFRX1 \block_r_reg[0][71]  ( .D(n3705), .CK(clk), .RN(n4241), .QN(n1017) );
  DFFRX1 \block_r_reg[6][71]  ( .D(n2937), .CK(clk), .RN(n4241), .QN(n249) );
  DFFRX1 \block_r_reg[4][71]  ( .D(n3193), .CK(clk), .RN(n4241), .QN(n505) );
  DFFRX1 \block_r_reg[2][71]  ( .D(n3449), .CK(clk), .RN(n4241), .QN(n761) );
  DFFRX1 \block_r_reg[0][70]  ( .D(n3706), .CK(clk), .RN(n4241), .QN(n1018) );
  DFFRX1 \block_r_reg[6][70]  ( .D(n2938), .CK(clk), .RN(n4241), .QN(n250) );
  DFFRX1 \block_r_reg[4][70]  ( .D(n3194), .CK(clk), .RN(n4240), .QN(n506) );
  DFFRX1 \block_r_reg[2][70]  ( .D(n3450), .CK(clk), .RN(n4240), .QN(n762) );
  DFFRX1 \block_r_reg[0][69]  ( .D(n3707), .CK(clk), .RN(n4240), .QN(n1019) );
  DFFRX1 \block_r_reg[6][69]  ( .D(n2939), .CK(clk), .RN(n4240), .QN(n251) );
  DFFRX1 \block_r_reg[4][69]  ( .D(n3195), .CK(clk), .RN(n4240), .QN(n507) );
  DFFRX1 \block_r_reg[2][69]  ( .D(n3451), .CK(clk), .RN(n4240), .QN(n763) );
  DFFRX1 \block_r_reg[0][68]  ( .D(n3708), .CK(clk), .RN(n4239), .QN(n1020) );
  DFFRX1 \block_r_reg[6][68]  ( .D(n2940), .CK(clk), .RN(n4239), .QN(n252) );
  DFFRX1 \block_r_reg[4][68]  ( .D(n3196), .CK(clk), .RN(n4239), .QN(n508) );
  DFFRX1 \block_r_reg[2][68]  ( .D(n3452), .CK(clk), .RN(n4239), .QN(n764) );
  DFFRX1 \block_r_reg[0][67]  ( .D(n3709), .CK(clk), .RN(n4239), .QN(n1021) );
  DFFRX1 \block_r_reg[6][67]  ( .D(n2941), .CK(clk), .RN(n4239), .QN(n253) );
  DFFRX1 \block_r_reg[4][67]  ( .D(n3197), .CK(clk), .RN(n4238), .QN(n509) );
  DFFRX1 \block_r_reg[2][67]  ( .D(n3453), .CK(clk), .RN(n4238), .QN(n765) );
  DFFRX1 \block_r_reg[0][66]  ( .D(n3710), .CK(clk), .RN(n4238), .QN(n1022) );
  DFFRX1 \block_r_reg[6][66]  ( .D(n2942), .CK(clk), .RN(n4238), .QN(n254) );
  DFFRX1 \block_r_reg[4][66]  ( .D(n3198), .CK(clk), .RN(n4238), .QN(n510) );
  DFFRX1 \block_r_reg[2][66]  ( .D(n3454), .CK(clk), .RN(n4238), .QN(n766) );
  DFFRX1 \block_r_reg[0][65]  ( .D(n3711), .CK(clk), .RN(n4237), .QN(n1023) );
  DFFRX1 \block_r_reg[6][65]  ( .D(n2943), .CK(clk), .RN(n4237), .QN(n255) );
  DFFRX1 \block_r_reg[4][65]  ( .D(n3199), .CK(clk), .RN(n4237), .QN(n511) );
  DFFRX1 \block_r_reg[2][65]  ( .D(n3455), .CK(clk), .RN(n4237), .QN(n767) );
  DFFRX1 \block_r_reg[0][64]  ( .D(n3712), .CK(clk), .RN(n4237), .QN(n1024) );
  DFFRX1 \block_r_reg[6][64]  ( .D(n2944), .CK(clk), .RN(n4237), .QN(n256) );
  DFFRX1 \block_r_reg[4][64]  ( .D(n3200), .CK(clk), .RN(n4236), .QN(n512) );
  DFFRX1 \block_r_reg[2][64]  ( .D(n3456), .CK(clk), .RN(n4236), .QN(n768) );
  DFFRX1 \block_r_reg[0][63]  ( .D(n3713), .CK(clk), .RN(n4236), .QN(n1025) );
  DFFRX1 \block_r_reg[6][63]  ( .D(n2945), .CK(clk), .RN(n4236), .QN(n257) );
  DFFRX1 \block_r_reg[4][63]  ( .D(n3201), .CK(clk), .RN(n4236), .QN(n513) );
  DFFRX1 \block_r_reg[2][63]  ( .D(n3457), .CK(clk), .RN(n4236), .QN(n769) );
  DFFRX1 \block_r_reg[0][62]  ( .D(n3714), .CK(clk), .RN(n4235), .QN(n1026) );
  DFFRX1 \block_r_reg[6][62]  ( .D(n2946), .CK(clk), .RN(n4235), .QN(n258) );
  DFFRX1 \block_r_reg[4][62]  ( .D(n3202), .CK(clk), .RN(n4235), .QN(n514) );
  DFFRX1 \block_r_reg[2][62]  ( .D(n3458), .CK(clk), .RN(n4235), .QN(n770) );
  DFFRX1 \block_r_reg[0][61]  ( .D(n3715), .CK(clk), .RN(n4235), .QN(n1027) );
  DFFRX1 \block_r_reg[6][61]  ( .D(n2947), .CK(clk), .RN(n4235), .QN(n259) );
  DFFRX1 \block_r_reg[4][61]  ( .D(n3203), .CK(clk), .RN(n4234), .QN(n515) );
  DFFRX1 \block_r_reg[2][61]  ( .D(n3459), .CK(clk), .RN(n4234), .QN(n771) );
  DFFRX1 \block_r_reg[0][60]  ( .D(n3716), .CK(clk), .RN(n4234), .QN(n1028) );
  DFFRX1 \block_r_reg[6][60]  ( .D(n2948), .CK(clk), .RN(n4234), .QN(n260) );
  DFFRX1 \block_r_reg[4][60]  ( .D(n3204), .CK(clk), .RN(n4234), .QN(n516) );
  DFFRX1 \block_r_reg[2][60]  ( .D(n3460), .CK(clk), .RN(n4234), .QN(n772) );
  DFFRX1 \block_r_reg[0][59]  ( .D(n3717), .CK(clk), .RN(n4233), .QN(n1029) );
  DFFRX1 \block_r_reg[6][59]  ( .D(n2949), .CK(clk), .RN(n4233), .QN(n261) );
  DFFRX1 \block_r_reg[4][59]  ( .D(n3205), .CK(clk), .RN(n4233), .QN(n517) );
  DFFRX1 \block_r_reg[2][59]  ( .D(n3461), .CK(clk), .RN(n4233), .QN(n773) );
  DFFRX1 \block_r_reg[0][58]  ( .D(n3718), .CK(clk), .RN(n4233), .QN(n1030) );
  DFFRX1 \block_r_reg[6][58]  ( .D(n2950), .CK(clk), .RN(n4233), .QN(n262) );
  DFFRX1 \block_r_reg[4][58]  ( .D(n3206), .CK(clk), .RN(n4232), .QN(n518) );
  DFFRX1 \block_r_reg[2][58]  ( .D(n3462), .CK(clk), .RN(n4232), .QN(n774) );
  DFFRX1 \block_r_reg[0][57]  ( .D(n3719), .CK(clk), .RN(n4232), .QN(n1031) );
  DFFRX1 \block_r_reg[6][57]  ( .D(n2951), .CK(clk), .RN(n4232), .QN(n263) );
  DFFRX1 \block_r_reg[4][57]  ( .D(n3207), .CK(clk), .RN(n4232), .QN(n519) );
  DFFRX1 \block_r_reg[2][57]  ( .D(n3463), .CK(clk), .RN(n4232), .QN(n775) );
  DFFRX1 \block_r_reg[0][56]  ( .D(n3720), .CK(clk), .RN(n4231), .QN(n1032) );
  DFFRX1 \block_r_reg[6][56]  ( .D(n2952), .CK(clk), .RN(n4231), .QN(n264) );
  DFFRX1 \block_r_reg[4][56]  ( .D(n3208), .CK(clk), .RN(n4231), .QN(n520) );
  DFFRX1 \block_r_reg[2][56]  ( .D(n3464), .CK(clk), .RN(n4231), .QN(n776) );
  DFFRX1 \block_r_reg[0][55]  ( .D(n3721), .CK(clk), .RN(n4231), .QN(n1033) );
  DFFRX1 \block_r_reg[6][55]  ( .D(n2953), .CK(clk), .RN(n4231), .QN(n265) );
  DFFRX1 \block_r_reg[4][55]  ( .D(n3209), .CK(clk), .RN(n4230), .QN(n521) );
  DFFRX1 \block_r_reg[2][55]  ( .D(n3465), .CK(clk), .RN(n4230), .QN(n777) );
  DFFRX1 \block_r_reg[0][54]  ( .D(n3722), .CK(clk), .RN(n4230), .QN(n1034) );
  DFFRX1 \block_r_reg[6][54]  ( .D(n2954), .CK(clk), .RN(n4230), .QN(n266) );
  DFFRX1 \block_r_reg[4][54]  ( .D(n3210), .CK(clk), .RN(n4230), .QN(n522) );
  DFFRX1 \block_r_reg[2][54]  ( .D(n3466), .CK(clk), .RN(n4230), .QN(n778) );
  DFFRX1 \block_r_reg[0][53]  ( .D(n3723), .CK(clk), .RN(n4229), .QN(n1035) );
  DFFRX1 \block_r_reg[6][53]  ( .D(n2955), .CK(clk), .RN(n4229), .QN(n267) );
  DFFRX1 \block_r_reg[4][53]  ( .D(n3211), .CK(clk), .RN(n4229), .QN(n523) );
  DFFRX1 \block_r_reg[2][53]  ( .D(n3467), .CK(clk), .RN(n4229), .QN(n779) );
  DFFRX1 \block_r_reg[0][52]  ( .D(n3724), .CK(clk), .RN(n4229), .QN(n1036) );
  DFFRX1 \block_r_reg[6][52]  ( .D(n2956), .CK(clk), .RN(n4229), .QN(n268) );
  DFFRX1 \block_r_reg[4][52]  ( .D(n3212), .CK(clk), .RN(n4228), .QN(n524) );
  DFFRX1 \block_r_reg[2][52]  ( .D(n3468), .CK(clk), .RN(n4228), .QN(n780) );
  DFFRX1 \block_r_reg[0][51]  ( .D(n3725), .CK(clk), .RN(n4228), .QN(n1037) );
  DFFRX1 \block_r_reg[6][51]  ( .D(n2957), .CK(clk), .RN(n4228), .QN(n269) );
  DFFRX1 \block_r_reg[4][51]  ( .D(n3213), .CK(clk), .RN(n4228), .QN(n525) );
  DFFRX1 \block_r_reg[2][51]  ( .D(n3469), .CK(clk), .RN(n4228), .QN(n781) );
  DFFRX1 \block_r_reg[0][50]  ( .D(n3726), .CK(clk), .RN(n4227), .QN(n1038) );
  DFFRX1 \block_r_reg[6][50]  ( .D(n2958), .CK(clk), .RN(n4227), .QN(n270) );
  DFFRX1 \block_r_reg[4][50]  ( .D(n3214), .CK(clk), .RN(n4227), .QN(n526) );
  DFFRX1 \block_r_reg[2][50]  ( .D(n3470), .CK(clk), .RN(n4227), .QN(n782) );
  DFFRX1 \block_r_reg[0][49]  ( .D(n3727), .CK(clk), .RN(n4227), .QN(n1039) );
  DFFRX1 \block_r_reg[6][49]  ( .D(n2959), .CK(clk), .RN(n4227), .QN(n271) );
  DFFRX1 \block_r_reg[4][49]  ( .D(n3215), .CK(clk), .RN(n4226), .QN(n527) );
  DFFRX1 \block_r_reg[2][49]  ( .D(n3471), .CK(clk), .RN(n4226), .QN(n783) );
  DFFRX1 \block_r_reg[0][48]  ( .D(n3728), .CK(clk), .RN(n4226), .QN(n1040) );
  DFFRX1 \block_r_reg[6][48]  ( .D(n2960), .CK(clk), .RN(n4226), .QN(n272) );
  DFFRX1 \block_r_reg[4][48]  ( .D(n3216), .CK(clk), .RN(n4226), .QN(n528) );
  DFFRX1 \block_r_reg[2][48]  ( .D(n3472), .CK(clk), .RN(n4226), .QN(n784) );
  DFFRX1 \block_r_reg[0][47]  ( .D(n3729), .CK(clk), .RN(n4225), .QN(n1041) );
  DFFRX1 \block_r_reg[6][47]  ( .D(n2961), .CK(clk), .RN(n4225), .QN(n273) );
  DFFRX1 \block_r_reg[4][47]  ( .D(n3217), .CK(clk), .RN(n4225), .QN(n529) );
  DFFRX1 \block_r_reg[2][47]  ( .D(n3473), .CK(clk), .RN(n4225), .QN(n785) );
  DFFRX1 \block_r_reg[0][46]  ( .D(n3730), .CK(clk), .RN(n4225), .QN(n1042) );
  DFFRX1 \block_r_reg[6][46]  ( .D(n2962), .CK(clk), .RN(n4225), .QN(n274) );
  DFFRX1 \block_r_reg[4][46]  ( .D(n3218), .CK(clk), .RN(n4224), .QN(n530) );
  DFFRX1 \block_r_reg[2][46]  ( .D(n3474), .CK(clk), .RN(n4224), .QN(n786) );
  DFFRX1 \block_r_reg[0][45]  ( .D(n3731), .CK(clk), .RN(n4224), .QN(n1043) );
  DFFRX1 \block_r_reg[6][45]  ( .D(n2963), .CK(clk), .RN(n4224), .QN(n275) );
  DFFRX1 \block_r_reg[4][45]  ( .D(n3219), .CK(clk), .RN(n4224), .QN(n531) );
  DFFRX1 \block_r_reg[2][45]  ( .D(n3475), .CK(clk), .RN(n4224), .QN(n787) );
  DFFRX1 \block_r_reg[0][44]  ( .D(n3732), .CK(clk), .RN(n4223), .QN(n1044) );
  DFFRX1 \block_r_reg[6][44]  ( .D(n2964), .CK(clk), .RN(n4223), .QN(n276) );
  DFFRX1 \block_r_reg[4][44]  ( .D(n3220), .CK(clk), .RN(n4223), .QN(n532) );
  DFFRX1 \block_r_reg[2][44]  ( .D(n3476), .CK(clk), .RN(n4223), .QN(n788) );
  DFFRX1 \block_r_reg[0][43]  ( .D(n3733), .CK(clk), .RN(n4223), .QN(n1045) );
  DFFRX1 \block_r_reg[6][43]  ( .D(n2965), .CK(clk), .RN(n4223), .QN(n277) );
  DFFRX1 \block_r_reg[4][43]  ( .D(n3221), .CK(clk), .RN(n4222), .QN(n533) );
  DFFRX1 \block_r_reg[2][43]  ( .D(n3477), .CK(clk), .RN(n4222), .QN(n789) );
  DFFRX1 \block_r_reg[0][42]  ( .D(n3734), .CK(clk), .RN(n4222), .QN(n1046) );
  DFFRX1 \block_r_reg[6][42]  ( .D(n2966), .CK(clk), .RN(n4222), .QN(n278) );
  DFFRX1 \block_r_reg[4][42]  ( .D(n3222), .CK(clk), .RN(n4222), .QN(n534) );
  DFFRX1 \block_r_reg[2][42]  ( .D(n3478), .CK(clk), .RN(n4222), .QN(n790) );
  DFFRX1 \block_r_reg[0][41]  ( .D(n3735), .CK(clk), .RN(n4221), .QN(n1047) );
  DFFRX1 \block_r_reg[6][41]  ( .D(n2967), .CK(clk), .RN(n4221), .QN(n279) );
  DFFRX1 \block_r_reg[4][41]  ( .D(n3223), .CK(clk), .RN(n4221), .QN(n535) );
  DFFRX1 \block_r_reg[2][41]  ( .D(n3479), .CK(clk), .RN(n4221), .QN(n791) );
  DFFRX1 \block_r_reg[0][40]  ( .D(n3736), .CK(clk), .RN(n4221), .QN(n1048) );
  DFFRX1 \block_r_reg[6][40]  ( .D(n2968), .CK(clk), .RN(n4221), .QN(n280) );
  DFFRX1 \block_r_reg[4][40]  ( .D(n3224), .CK(clk), .RN(n4220), .QN(n536) );
  DFFRX1 \block_r_reg[2][40]  ( .D(n3480), .CK(clk), .RN(n4220), .QN(n792) );
  DFFRX1 \block_r_reg[0][39]  ( .D(n3737), .CK(clk), .RN(n4220), .QN(n1049) );
  DFFRX1 \block_r_reg[6][39]  ( .D(n2969), .CK(clk), .RN(n4220), .QN(n281) );
  DFFRX1 \block_r_reg[4][39]  ( .D(n3225), .CK(clk), .RN(n4220), .QN(n537) );
  DFFRX1 \block_r_reg[2][39]  ( .D(n3481), .CK(clk), .RN(n4220), .QN(n793) );
  DFFRX1 \block_r_reg[0][38]  ( .D(n3738), .CK(clk), .RN(n4219), .QN(n1050) );
  DFFRX1 \block_r_reg[6][38]  ( .D(n2970), .CK(clk), .RN(n4219), .QN(n282) );
  DFFRX1 \block_r_reg[4][38]  ( .D(n3226), .CK(clk), .RN(n4219), .QN(n538) );
  DFFRX1 \block_r_reg[2][38]  ( .D(n3482), .CK(clk), .RN(n4219), .QN(n794) );
  DFFRX1 \block_r_reg[0][37]  ( .D(n3739), .CK(clk), .RN(n4219), .QN(n1051) );
  DFFRX1 \block_r_reg[6][37]  ( .D(n2971), .CK(clk), .RN(n4219), .QN(n283) );
  DFFRX1 \block_r_reg[4][37]  ( .D(n3227), .CK(clk), .RN(n4218), .QN(n539) );
  DFFRX1 \block_r_reg[2][37]  ( .D(n3483), .CK(clk), .RN(n4218), .QN(n795) );
  DFFRX1 \block_r_reg[0][36]  ( .D(n3740), .CK(clk), .RN(n4218), .QN(n1052) );
  DFFRX1 \block_r_reg[6][36]  ( .D(n2972), .CK(clk), .RN(n4218), .QN(n284) );
  DFFRX1 \block_r_reg[4][36]  ( .D(n3228), .CK(clk), .RN(n4218), .QN(n540) );
  DFFRX1 \block_r_reg[2][36]  ( .D(n3484), .CK(clk), .RN(n4218), .QN(n796) );
  DFFRX1 \block_r_reg[0][35]  ( .D(n3741), .CK(clk), .RN(n4217), .QN(n1053) );
  DFFRX1 \block_r_reg[6][35]  ( .D(n2973), .CK(clk), .RN(n4217), .QN(n285) );
  DFFRX1 \block_r_reg[4][35]  ( .D(n3229), .CK(clk), .RN(n4217), .QN(n541) );
  DFFRX1 \block_r_reg[2][35]  ( .D(n3485), .CK(clk), .RN(n4217), .QN(n797) );
  DFFRX1 \block_r_reg[0][34]  ( .D(n3742), .CK(clk), .RN(n4217), .QN(n1054) );
  DFFRX1 \block_r_reg[6][34]  ( .D(n2974), .CK(clk), .RN(n4217), .QN(n286) );
  DFFRX1 \block_r_reg[2][34]  ( .D(n3486), .CK(clk), .RN(n4216), .QN(n798) );
  DFFRX1 \block_r_reg[0][33]  ( .D(n3743), .CK(clk), .RN(n4216), .QN(n1055) );
  DFFRX1 \block_r_reg[6][33]  ( .D(n2975), .CK(clk), .RN(n4216), .QN(n287) );
  DFFRX1 \block_r_reg[2][33]  ( .D(n3487), .CK(clk), .RN(n4216), .QN(n799) );
  DFFRX1 \block_r_reg[0][32]  ( .D(n3744), .CK(clk), .RN(n4215), .QN(n1056) );
  DFFRX1 \block_r_reg[6][32]  ( .D(n2976), .CK(clk), .RN(n4215), .QN(n288) );
  DFFRX1 \block_r_reg[2][32]  ( .D(n3488), .CK(clk), .RN(n4215), .QN(n800) );
  DFFRX1 \block_r_reg[0][31]  ( .D(n3745), .CK(clk), .RN(n4215), .QN(n1057) );
  DFFRX1 \block_r_reg[6][31]  ( .D(n2977), .CK(clk), .RN(n4215), .QN(n289) );
  DFFRX1 \block_r_reg[2][31]  ( .D(n3489), .CK(clk), .RN(n4214), .QN(n801) );
  DFFRX1 \block_r_reg[0][30]  ( .D(n3746), .CK(clk), .RN(n4214), .QN(n1058) );
  DFFRX1 \block_r_reg[6][30]  ( .D(n2978), .CK(clk), .RN(n4214), .QN(n290) );
  DFFRX1 \block_r_reg[2][30]  ( .D(n3490), .CK(clk), .RN(n4214), .QN(n802) );
  DFFRX1 \block_r_reg[0][29]  ( .D(n3747), .CK(clk), .RN(n4213), .QN(n1059) );
  DFFRX1 \block_r_reg[6][29]  ( .D(n2979), .CK(clk), .RN(n4213), .QN(n291) );
  DFFRX1 \block_r_reg[2][29]  ( .D(n3491), .CK(clk), .RN(n4213), .QN(n803) );
  DFFRX1 \block_r_reg[0][28]  ( .D(n3748), .CK(clk), .RN(n4213), .QN(n1060) );
  DFFRX1 \block_r_reg[6][28]  ( .D(n2980), .CK(clk), .RN(n4213), .QN(n292) );
  DFFRX1 \block_r_reg[2][28]  ( .D(n3492), .CK(clk), .RN(n4212), .QN(n804) );
  DFFRX1 \block_r_reg[0][27]  ( .D(n3749), .CK(clk), .RN(n4212), .QN(n1061) );
  DFFRX1 \block_r_reg[6][27]  ( .D(n2981), .CK(clk), .RN(n4212), .QN(n293) );
  DFFRX1 \block_r_reg[2][27]  ( .D(n3493), .CK(clk), .RN(n4212), .QN(n805) );
  DFFRX1 \block_r_reg[0][26]  ( .D(n3750), .CK(clk), .RN(n4211), .QN(n1062) );
  DFFRX1 \block_r_reg[6][26]  ( .D(n2982), .CK(clk), .RN(n4211), .QN(n294) );
  DFFRX1 \block_r_reg[2][26]  ( .D(n3494), .CK(clk), .RN(n4211), .QN(n806) );
  DFFRX1 \block_r_reg[0][25]  ( .D(n3751), .CK(clk), .RN(n4211), .QN(n1063) );
  DFFRX1 \block_r_reg[6][25]  ( .D(n2983), .CK(clk), .RN(n4211), .QN(n295) );
  DFFRX1 \block_r_reg[2][25]  ( .D(n3495), .CK(clk), .RN(n4210), .QN(n807) );
  DFFRX1 \block_r_reg[0][24]  ( .D(n3752), .CK(clk), .RN(n4210), .QN(n1064) );
  DFFRX1 \block_r_reg[6][24]  ( .D(n2984), .CK(clk), .RN(n4210), .QN(n296) );
  DFFRX1 \block_r_reg[2][24]  ( .D(n3496), .CK(clk), .RN(n4210), .QN(n808) );
  DFFRX1 \block_r_reg[0][23]  ( .D(n3753), .CK(clk), .RN(n4209), .QN(n1065) );
  DFFRX1 \block_r_reg[6][23]  ( .D(n2985), .CK(clk), .RN(n4209), .QN(n297) );
  DFFRX1 \block_r_reg[2][23]  ( .D(n3497), .CK(clk), .RN(n4209), .QN(n809) );
  DFFRX1 \block_r_reg[0][22]  ( .D(n3754), .CK(clk), .RN(n4209), .QN(n1066) );
  DFFRX1 \block_r_reg[6][22]  ( .D(n2986), .CK(clk), .RN(n4209), .QN(n298) );
  DFFRX1 \block_r_reg[2][22]  ( .D(n3498), .CK(clk), .RN(n4208), .QN(n810) );
  DFFRX1 \block_r_reg[0][21]  ( .D(n3755), .CK(clk), .RN(n4208), .QN(n1067) );
  DFFRX1 \block_r_reg[6][21]  ( .D(n2987), .CK(clk), .RN(n4208), .QN(n299) );
  DFFRX1 \block_r_reg[2][21]  ( .D(n3499), .CK(clk), .RN(n4208), .QN(n811) );
  DFFRX1 \block_r_reg[0][20]  ( .D(n3756), .CK(clk), .RN(n4207), .QN(n1068) );
  DFFRX1 \block_r_reg[6][20]  ( .D(n2988), .CK(clk), .RN(n4207), .QN(n300) );
  DFFRX1 \block_r_reg[2][20]  ( .D(n3500), .CK(clk), .RN(n4207), .QN(n812) );
  DFFRX1 \block_r_reg[0][19]  ( .D(n3757), .CK(clk), .RN(n4207), .QN(n1069) );
  DFFRX1 \block_r_reg[6][19]  ( .D(n2989), .CK(clk), .RN(n4207), .QN(n301) );
  DFFRX1 \block_r_reg[2][19]  ( .D(n3501), .CK(clk), .RN(n4206), .QN(n813) );
  DFFRX1 \block_r_reg[0][18]  ( .D(n3758), .CK(clk), .RN(n4206), .QN(n1070) );
  DFFRX1 \block_r_reg[6][18]  ( .D(n2990), .CK(clk), .RN(n4206), .QN(n302) );
  DFFRX1 \block_r_reg[4][18]  ( .D(n3246), .CK(clk), .RN(n4206), .QN(n558) );
  DFFRX1 \block_r_reg[2][18]  ( .D(n3502), .CK(clk), .RN(n4206), .QN(n814) );
  DFFRX1 \tag_r_reg[0][0]  ( .D(n3994), .CK(clk), .RN(n4309), .Q(\tag_r[0][0] ), .QN(n1288) );
  DFFRX1 \tag_r_reg[1][18]  ( .D(n3807), .CK(clk), .RN(n4307), .Q(
        \tag_r[1][18] ), .QN(n1245) );
  DFFRX1 \tag_r_reg[1][17]  ( .D(n3808), .CK(clk), .RN(n4307), .Q(
        \tag_r[1][17] ), .QN(n1246) );
  DFFRX1 \tag_r_reg[1][16]  ( .D(n3809), .CK(clk), .RN(n4307), .Q(
        \tag_r[1][16] ), .QN(n1247) );
  DFFRX1 \tag_r_reg[1][15]  ( .D(n3810), .CK(clk), .RN(n4307), .Q(
        \tag_r[1][15] ), .QN(n1248) );
  DFFRX1 \tag_r_reg[1][14]  ( .D(n3811), .CK(clk), .RN(n4307), .Q(
        \tag_r[1][14] ), .QN(n1249) );
  DFFRX1 \tag_r_reg[1][13]  ( .D(n3812), .CK(clk), .RN(n4306), .Q(
        \tag_r[1][13] ), .QN(n1250) );
  DFFRX1 \tag_r_reg[1][12]  ( .D(n3813), .CK(clk), .RN(n4306), .Q(
        \tag_r[1][12] ), .QN(n1251) );
  DFFRX1 \tag_r_reg[1][6]  ( .D(n3819), .CK(clk), .RN(n4306), .Q(\tag_r[1][6] ), .QN(n1257) );
  DFFRX1 \tag_r_reg[1][4]  ( .D(n3821), .CK(clk), .RN(n4306), .Q(\tag_r[1][4] ), .QN(n1259) );
  DFFRX1 \tag_r_reg[1][3]  ( .D(n3822), .CK(clk), .RN(n4306), .Q(\tag_r[1][3] ), .QN(n1260) );
  DFFRX1 \tag_r_reg[1][2]  ( .D(n3823), .CK(clk), .RN(n4306), .Q(\tag_r[1][2] ), .QN(n1261) );
  DFFRX1 \tag_r_reg[1][1]  ( .D(n3824), .CK(clk), .RN(n4305), .Q(\tag_r[1][1] ), .QN(n1262) );
  DFFRX1 \tag_r_reg[1][0]  ( .D(n3825), .CK(clk), .RN(n4305), .Q(\tag_r[1][0] ), .QN(n1263) );
  DFFRX1 \tag_r_reg[2][18]  ( .D(n3832), .CK(clk), .RN(n4305), .Q(
        \tag_r[2][18] ), .QN(n1220) );
  DFFRX1 \tag_r_reg[2][17]  ( .D(n3833), .CK(clk), .RN(n4305), .Q(
        \tag_r[2][17] ), .QN(n1221) );
  DFFRX1 \tag_r_reg[2][16]  ( .D(n3834), .CK(clk), .RN(n4305), .Q(
        \tag_r[2][16] ), .QN(n1222) );
  DFFRX1 \tag_r_reg[2][15]  ( .D(n3835), .CK(clk), .RN(n4305), .Q(
        \tag_r[2][15] ), .QN(n1223) );
  DFFRX1 \tag_r_reg[2][14]  ( .D(n3836), .CK(clk), .RN(n4304), .Q(
        \tag_r[2][14] ), .QN(n1224) );
  DFFRX1 \tag_r_reg[2][13]  ( .D(n3837), .CK(clk), .RN(n4304), .Q(
        \tag_r[2][13] ), .QN(n1225) );
  DFFRX1 \tag_r_reg[2][12]  ( .D(n3838), .CK(clk), .RN(n4304), .Q(
        \tag_r[2][12] ), .QN(n1226) );
  DFFRX1 \tag_r_reg[2][6]  ( .D(n3844), .CK(clk), .RN(n4304), .Q(\tag_r[2][6] ), .QN(n1232) );
  DFFRX1 \tag_r_reg[2][4]  ( .D(n3846), .CK(clk), .RN(n4304), .Q(\tag_r[2][4] ), .QN(n1234) );
  DFFRX1 \tag_r_reg[2][3]  ( .D(n3847), .CK(clk), .RN(n4304), .Q(\tag_r[2][3] ), .QN(n1235) );
  DFFRX1 \tag_r_reg[2][2]  ( .D(n3848), .CK(clk), .RN(n4303), .Q(\tag_r[2][2] ), .QN(n1236) );
  DFFRX1 \tag_r_reg[2][1]  ( .D(n3849), .CK(clk), .RN(n4303), .Q(\tag_r[2][1] ), .QN(n1237) );
  DFFRX1 \tag_r_reg[2][0]  ( .D(n3850), .CK(clk), .RN(n4303), .Q(\tag_r[2][0] ), .QN(n1238) );
  DFFRX1 \tag_r_reg[3][18]  ( .D(n3857), .CK(clk), .RN(n4303), .Q(
        \tag_r[3][18] ), .QN(n1195) );
  DFFRX1 \tag_r_reg[3][17]  ( .D(n3858), .CK(clk), .RN(n4303), .Q(
        \tag_r[3][17] ), .QN(n1196) );
  DFFRX1 \tag_r_reg[3][16]  ( .D(n3859), .CK(clk), .RN(n4303), .Q(
        \tag_r[3][16] ), .QN(n1197) );
  DFFRX1 \tag_r_reg[3][15]  ( .D(n3860), .CK(clk), .RN(n4302), .Q(
        \tag_r[3][15] ), .QN(n1198) );
  DFFRX1 \tag_r_reg[3][14]  ( .D(n3861), .CK(clk), .RN(n4302), .Q(
        \tag_r[3][14] ), .QN(n1199) );
  DFFRX1 \tag_r_reg[3][13]  ( .D(n3862), .CK(clk), .RN(n4302), .Q(
        \tag_r[3][13] ), .QN(n1200) );
  DFFRX1 \tag_r_reg[3][12]  ( .D(n3863), .CK(clk), .RN(n4302), .Q(
        \tag_r[3][12] ), .QN(n1201) );
  DFFRX1 \tag_r_reg[3][6]  ( .D(n3869), .CK(clk), .RN(n4302), .Q(\tag_r[3][6] ), .QN(n1207) );
  DFFRX1 \tag_r_reg[3][4]  ( .D(n3871), .CK(clk), .RN(n4302), .Q(\tag_r[3][4] ), .QN(n1209) );
  DFFRX1 \tag_r_reg[3][3]  ( .D(n3872), .CK(clk), .RN(n4301), .Q(\tag_r[3][3] ), .QN(n1210) );
  DFFRX1 \tag_r_reg[3][2]  ( .D(n3873), .CK(clk), .RN(n4301), .Q(\tag_r[3][2] ), .QN(n1211) );
  DFFRX1 \tag_r_reg[3][1]  ( .D(n3874), .CK(clk), .RN(n4301), .Q(\tag_r[3][1] ), .QN(n1212) );
  DFFRX1 \tag_r_reg[3][0]  ( .D(n3875), .CK(clk), .RN(n4301), .Q(\tag_r[3][0] ), .QN(n1213) );
  DFFRX1 \tag_r_reg[4][18]  ( .D(n3882), .CK(clk), .RN(n4301), .Q(
        \tag_r[4][18] ), .QN(n1170) );
  DFFRX1 \tag_r_reg[4][17]  ( .D(n3883), .CK(clk), .RN(n4301), .Q(
        \tag_r[4][17] ), .QN(n1171) );
  DFFRX1 \tag_r_reg[4][16]  ( .D(n3884), .CK(clk), .RN(n4300), .Q(
        \tag_r[4][16] ), .QN(n1172) );
  DFFRX1 \tag_r_reg[4][15]  ( .D(n3885), .CK(clk), .RN(n4300), .Q(
        \tag_r[4][15] ), .QN(n1173) );
  DFFRX1 \tag_r_reg[4][14]  ( .D(n3886), .CK(clk), .RN(n4300), .Q(
        \tag_r[4][14] ), .QN(n1174) );
  DFFRX1 \tag_r_reg[4][13]  ( .D(n3887), .CK(clk), .RN(n4300), .Q(
        \tag_r[4][13] ), .QN(n1175) );
  DFFRX1 \tag_r_reg[4][12]  ( .D(n3888), .CK(clk), .RN(n4300), .Q(
        \tag_r[4][12] ), .QN(n1176) );
  DFFRX1 \tag_r_reg[4][6]  ( .D(n3894), .CK(clk), .RN(n4300), .Q(\tag_r[4][6] ), .QN(n1182) );
  DFFRX1 \tag_r_reg[4][4]  ( .D(n3896), .CK(clk), .RN(n4299), .Q(\tag_r[4][4] ), .QN(n1184) );
  DFFRX1 \tag_r_reg[4][3]  ( .D(n3897), .CK(clk), .RN(n4299), .Q(\tag_r[4][3] ), .QN(n1185) );
  DFFRX1 \tag_r_reg[4][2]  ( .D(n3898), .CK(clk), .RN(n4299), .Q(\tag_r[4][2] ), .QN(n1186) );
  DFFRX1 \tag_r_reg[4][1]  ( .D(n3899), .CK(clk), .RN(n4299), .Q(\tag_r[4][1] ), .QN(n1187) );
  DFFRX1 \tag_r_reg[4][0]  ( .D(n3900), .CK(clk), .RN(n4299), .Q(\tag_r[4][0] ), .QN(n1188) );
  DFFRX1 \tag_r_reg[5][18]  ( .D(n3907), .CK(clk), .RN(n4299), .Q(
        \tag_r[5][18] ), .QN(n1145) );
  DFFRX1 \tag_r_reg[5][17]  ( .D(n3908), .CK(clk), .RN(n4298), .Q(
        \tag_r[5][17] ), .QN(n1146) );
  DFFRX1 \tag_r_reg[5][16]  ( .D(n3909), .CK(clk), .RN(n4298), .Q(
        \tag_r[5][16] ), .QN(n1147) );
  DFFRX1 \tag_r_reg[5][15]  ( .D(n3910), .CK(clk), .RN(n4298), .Q(
        \tag_r[5][15] ), .QN(n1148) );
  DFFRX1 \tag_r_reg[5][14]  ( .D(n3911), .CK(clk), .RN(n4298), .Q(
        \tag_r[5][14] ), .QN(n1149) );
  DFFRX1 \tag_r_reg[5][13]  ( .D(n3912), .CK(clk), .RN(n4298), .Q(
        \tag_r[5][13] ), .QN(n1150) );
  DFFRX1 \tag_r_reg[5][12]  ( .D(n3913), .CK(clk), .RN(n4298), .Q(
        \tag_r[5][12] ), .QN(n1151) );
  DFFRX1 \tag_r_reg[5][6]  ( .D(n3919), .CK(clk), .RN(n4298), .Q(\tag_r[5][6] ), .QN(n1157) );
  DFFRX1 \tag_r_reg[5][4]  ( .D(n3921), .CK(clk), .RN(n4297), .Q(\tag_r[5][4] ), .QN(n1159) );
  DFFRX1 \tag_r_reg[5][3]  ( .D(n3922), .CK(clk), .RN(n4297), .Q(\tag_r[5][3] ), .QN(n1160) );
  DFFRX1 \tag_r_reg[5][2]  ( .D(n3923), .CK(clk), .RN(n4297), .Q(\tag_r[5][2] ), .QN(n1161) );
  DFFRX1 \tag_r_reg[5][1]  ( .D(n3924), .CK(clk), .RN(n4297), .Q(\tag_r[5][1] ), .QN(n1162) );
  DFFRX1 \tag_r_reg[5][0]  ( .D(n3925), .CK(clk), .RN(n4297), .Q(\tag_r[5][0] ), .QN(n1163) );
  DFFRX1 \tag_r_reg[6][18]  ( .D(n3932), .CK(clk), .RN(n4296), .Q(
        \tag_r[6][18] ), .QN(n1120) );
  DFFRX1 \tag_r_reg[6][17]  ( .D(n3933), .CK(clk), .RN(n4296), .Q(
        \tag_r[6][17] ), .QN(n1121) );
  DFFRX1 \tag_r_reg[6][16]  ( .D(n3934), .CK(clk), .RN(n4296), .Q(
        \tag_r[6][16] ), .QN(n1122) );
  DFFRX1 \tag_r_reg[6][15]  ( .D(n3935), .CK(clk), .RN(n4296), .Q(
        \tag_r[6][15] ), .QN(n1123) );
  DFFRX1 \tag_r_reg[6][14]  ( .D(n3936), .CK(clk), .RN(n4296), .Q(
        \tag_r[6][14] ), .QN(n1124) );
  DFFRX1 \tag_r_reg[6][13]  ( .D(n3937), .CK(clk), .RN(n4296), .Q(
        \tag_r[6][13] ), .QN(n1125) );
  DFFRX1 \tag_r_reg[6][12]  ( .D(n3938), .CK(clk), .RN(n4296), .Q(
        \tag_r[6][12] ), .QN(n1126) );
  DFFRX1 \tag_r_reg[6][6]  ( .D(n3944), .CK(clk), .RN(n4295), .Q(\tag_r[6][6] ), .QN(n1132) );
  DFFRX1 \tag_r_reg[6][4]  ( .D(n3946), .CK(clk), .RN(n4295), .Q(\tag_r[6][4] ), .QN(n1134) );
  DFFRX1 \tag_r_reg[6][3]  ( .D(n3947), .CK(clk), .RN(n4295), .Q(\tag_r[6][3] ), .QN(n1135) );
  DFFRX1 \tag_r_reg[6][2]  ( .D(n3948), .CK(clk), .RN(n4295), .Q(\tag_r[6][2] ), .QN(n1136) );
  DFFRX1 \tag_r_reg[6][1]  ( .D(n3949), .CK(clk), .RN(n4295), .Q(\tag_r[6][1] ), .QN(n1137) );
  DFFRX1 \tag_r_reg[6][0]  ( .D(n3950), .CK(clk), .RN(n4295), .Q(\tag_r[6][0] ), .QN(n1138) );
  DFFRX1 \tag_r_reg[7][18]  ( .D(n3957), .CK(clk), .RN(n4294), .Q(
        \tag_r[7][18] ), .QN(n1095) );
  DFFRX1 \tag_r_reg[7][17]  ( .D(n3958), .CK(clk), .RN(n4294), .Q(
        \tag_r[7][17] ), .QN(n1096) );
  DFFRX1 \tag_r_reg[7][15]  ( .D(n3960), .CK(clk), .RN(n4294), .Q(
        \tag_r[7][15] ), .QN(n1098) );
  DFFRX1 \tag_r_reg[7][14]  ( .D(n3961), .CK(clk), .RN(n4294), .Q(
        \tag_r[7][14] ), .QN(n1099) );
  DFFRX1 \tag_r_reg[7][13]  ( .D(n3962), .CK(clk), .RN(n4294), .Q(
        \tag_r[7][13] ), .QN(n1100) );
  DFFRX1 \tag_r_reg[7][12]  ( .D(n3963), .CK(clk), .RN(n4294), .Q(
        \tag_r[7][12] ), .QN(n1101) );
  DFFRX1 \tag_r_reg[7][11]  ( .D(n3964), .CK(clk), .RN(n4294), .Q(
        \tag_r[7][11] ), .QN(n1102) );
  DFFRX1 \tag_r_reg[7][6]  ( .D(n3969), .CK(clk), .RN(n4293), .Q(\tag_r[7][6] ), .QN(n1107) );
  DFFRX1 \tag_r_reg[7][4]  ( .D(n3971), .CK(clk), .RN(n4293), .Q(\tag_r[7][4] ), .QN(n1109) );
  DFFRX1 \tag_r_reg[7][3]  ( .D(n3972), .CK(clk), .RN(n4293), .Q(\tag_r[7][3] ), .QN(n1110) );
  DFFRX1 \tag_r_reg[7][2]  ( .D(n3973), .CK(clk), .RN(n4293), .Q(\tag_r[7][2] ), .QN(n1111) );
  DFFRX1 \tag_r_reg[7][1]  ( .D(n3974), .CK(clk), .RN(n4293), .Q(\tag_r[7][1] ), .QN(n1112) );
  DFFRX1 \tag_r_reg[7][0]  ( .D(n3975), .CK(clk), .RN(n4293), .Q(\tag_r[7][0] ), .QN(n1113) );
  DFFRX1 \tag_r_reg[0][18]  ( .D(n3783), .CK(clk), .RN(n4292), .Q(
        \tag_r[0][18] ), .QN(n1270) );
  DFFRX1 \tag_r_reg[0][17]  ( .D(n3784), .CK(clk), .RN(n4292), .Q(
        \tag_r[0][17] ), .QN(n1271) );
  DFFRX1 \tag_r_reg[0][15]  ( .D(n3786), .CK(clk), .RN(n4292), .Q(
        \tag_r[0][15] ), .QN(n1273) );
  DFFRX1 \tag_r_reg[0][14]  ( .D(n3787), .CK(clk), .RN(n4292), .Q(
        \tag_r[0][14] ), .QN(n1274) );
  DFFRX1 \tag_r_reg[0][13]  ( .D(n3788), .CK(clk), .RN(n4292), .Q(
        \tag_r[0][13] ), .QN(n1275) );
  DFFRX1 \tag_r_reg[0][12]  ( .D(n3789), .CK(clk), .RN(n4292), .Q(
        \tag_r[0][12] ), .QN(n1276) );
  DFFRX1 \tag_r_reg[0][11]  ( .D(n3790), .CK(clk), .RN(n4292), .Q(
        \tag_r[0][11] ), .QN(n1277) );
  DFFRX1 \tag_r_reg[0][6]  ( .D(n3795), .CK(clk), .RN(n4291), .Q(\tag_r[0][6] ), .QN(n1282) );
  DFFRX1 \tag_r_reg[0][4]  ( .D(n3797), .CK(clk), .RN(n4291), .Q(\tag_r[0][4] ), .QN(n1284) );
  DFFRX1 \tag_r_reg[0][3]  ( .D(n3798), .CK(clk), .RN(n4291), .Q(\tag_r[0][3] ), .QN(n1285) );
  DFFRX1 \tag_r_reg[0][2]  ( .D(n3799), .CK(clk), .RN(n4291), .Q(\tag_r[0][2] ), .QN(n1286) );
  DFFRX1 \tag_r_reg[0][1]  ( .D(n3800), .CK(clk), .RN(n4291), .Q(\tag_r[0][1] ), .QN(n1287) );
  DFFRX1 \tag_r_reg[1][24]  ( .D(n3801), .CK(clk), .RN(n4307), .Q(n1306), .QN(
        n1239) );
  DFFRX1 \tag_r_reg[3][24]  ( .D(n3851), .CK(clk), .RN(n4303), .Q(n1304), .QN(
        n1189) );
  DFFRX1 \tag_r_reg[5][24]  ( .D(n3901), .CK(clk), .RN(n4299), .Q(n1302), .QN(
        n1139) );
  DFFRX1 \tag_r_reg[7][24]  ( .D(n3951), .CK(clk), .RN(n4295), .Q(n1301), .QN(
        n1089) );
  DFFRX1 \tag_r_reg[2][24]  ( .D(n3826), .CK(clk), .RN(n4305), .Q(n1305), .QN(
        n1214) );
  DFFRX1 \tag_r_reg[4][24]  ( .D(n3876), .CK(clk), .RN(n4301), .Q(n1303), .QN(
        n1164) );
  DFFRX1 \tag_r_reg[6][24]  ( .D(n3926), .CK(clk), .RN(n4297), .Q(n1307), .QN(
        n1114) );
  DFFRX1 \tag_r_reg[0][24]  ( .D(n3777), .CK(clk), .RN(n4293), .Q(n1300), .QN(
        n1264) );
  DFFRX1 \state_r_reg[0]  ( .D(n3992), .CK(clk), .RN(n4309), .Q(\state_r[0] ), 
        .QN(n64) );
  DFFRX1 \state_r_reg[1]  ( .D(n3993), .CK(clk), .RN(n4309), .Q(n4419), .QN(
        n61) );
  DFFRX1 \valid_r_reg[4]  ( .D(n3979), .CK(clk), .RN(n4308), .QN(n46) );
  DFFRX1 \dirty_r_reg[4]  ( .D(n3988), .CK(clk), .RN(n4308), .QN(n38) );
  DFFRX1 \valid_r_reg[6]  ( .D(n3977), .CK(clk), .RN(n4308), .QN(n44) );
  DFFRX1 \dirty_r_reg[6]  ( .D(n3990), .CK(clk), .RN(n4308), .QN(n36) );
  DFFRX1 \valid_r_reg[5]  ( .D(n3978), .CK(clk), .RN(n4308), .QN(n45) );
  DFFRX1 \dirty_r_reg[5]  ( .D(n3989), .CK(clk), .RN(n4308), .QN(n37) );
  DFFRX1 \valid_r_reg[7]  ( .D(n3976), .CK(clk), .RN(n4308), .QN(n43) );
  DFFRX1 \dirty_r_reg[7]  ( .D(n3991), .CK(clk), .RN(n4308), .QN(n35) );
  DFFRX1 \tag_r_reg[3][11]  ( .D(n3864), .CK(clk), .RN(n4302), .QN(n1202) );
  DFFRX1 \tag_r_reg[3][10]  ( .D(n3865), .CK(clk), .RN(n4302), .QN(n1203) );
  DFFRX1 \tag_r_reg[3][9]  ( .D(n3866), .CK(clk), .RN(n4302), .QN(n1204) );
  DFFRX1 \tag_r_reg[3][8]  ( .D(n3867), .CK(clk), .RN(n4302), .QN(n1205) );
  DFFRX1 \tag_r_reg[3][7]  ( .D(n3868), .CK(clk), .RN(n4302), .QN(n1206) );
  DFFRX1 \tag_r_reg[3][5]  ( .D(n3870), .CK(clk), .RN(n4302), .QN(n1208) );
  DFFRX1 \tag_r_reg[2][11]  ( .D(n3839), .CK(clk), .RN(n4304), .QN(n1227) );
  DFFRX1 \tag_r_reg[2][10]  ( .D(n3840), .CK(clk), .RN(n4304), .QN(n1228) );
  DFFRX1 \tag_r_reg[2][9]  ( .D(n3841), .CK(clk), .RN(n4304), .QN(n1229) );
  DFFRX1 \tag_r_reg[2][8]  ( .D(n3842), .CK(clk), .RN(n4304), .QN(n1230) );
  DFFRX1 \tag_r_reg[2][7]  ( .D(n3843), .CK(clk), .RN(n4304), .QN(n1231) );
  DFFRX1 \tag_r_reg[2][5]  ( .D(n3845), .CK(clk), .RN(n4304), .QN(n1233) );
  DFFRX1 \tag_r_reg[3][23]  ( .D(n3852), .CK(clk), .RN(n4303), .QN(n1190) );
  DFFRX1 \tag_r_reg[3][22]  ( .D(n3853), .CK(clk), .RN(n4303), .QN(n1191) );
  DFFRX1 \tag_r_reg[3][21]  ( .D(n3854), .CK(clk), .RN(n4303), .QN(n1192) );
  DFFRX1 \tag_r_reg[3][20]  ( .D(n3855), .CK(clk), .RN(n4303), .QN(n1193) );
  DFFRX1 \tag_r_reg[3][19]  ( .D(n3856), .CK(clk), .RN(n4303), .QN(n1194) );
  DFFRX1 \tag_r_reg[2][23]  ( .D(n3827), .CK(clk), .RN(n4305), .QN(n1215) );
  DFFRX1 \tag_r_reg[2][22]  ( .D(n3828), .CK(clk), .RN(n4305), .QN(n1216) );
  DFFRX1 \tag_r_reg[2][21]  ( .D(n3829), .CK(clk), .RN(n4305), .QN(n1217) );
  DFFRX1 \tag_r_reg[2][20]  ( .D(n3830), .CK(clk), .RN(n4305), .QN(n1218) );
  DFFRX1 \tag_r_reg[2][19]  ( .D(n3831), .CK(clk), .RN(n4305), .QN(n1219) );
  DFFRX1 \tag_r_reg[0][10]  ( .D(n3791), .CK(clk), .RN(n4292), .QN(n1278) );
  DFFRX1 \tag_r_reg[0][9]  ( .D(n3792), .CK(clk), .RN(n4292), .QN(n1279) );
  DFFRX1 \tag_r_reg[0][8]  ( .D(n3793), .CK(clk), .RN(n4291), .QN(n1280) );
  DFFRX1 \tag_r_reg[0][7]  ( .D(n3794), .CK(clk), .RN(n4291), .QN(n1281) );
  DFFRX1 \tag_r_reg[0][5]  ( .D(n3796), .CK(clk), .RN(n4291), .QN(n1283) );
  DFFRX1 \tag_r_reg[0][23]  ( .D(n3778), .CK(clk), .RN(n4293), .QN(n1265) );
  DFFRX1 \tag_r_reg[0][22]  ( .D(n3779), .CK(clk), .RN(n4293), .QN(n1266) );
  DFFRX1 \tag_r_reg[0][21]  ( .D(n3780), .CK(clk), .RN(n4293), .QN(n1267) );
  DFFRX1 \tag_r_reg[0][20]  ( .D(n3781), .CK(clk), .RN(n4292), .QN(n1268) );
  DFFRX1 \tag_r_reg[0][19]  ( .D(n3782), .CK(clk), .RN(n4292), .QN(n1269) );
  DFFRX1 \tag_r_reg[0][16]  ( .D(n3785), .CK(clk), .RN(n4292), .QN(n1272) );
  DFFRX1 \tag_r_reg[1][11]  ( .D(n3814), .CK(clk), .RN(n4306), .QN(n1252) );
  DFFRX1 \tag_r_reg[1][10]  ( .D(n3815), .CK(clk), .RN(n4306), .QN(n1253) );
  DFFRX1 \tag_r_reg[1][9]  ( .D(n3816), .CK(clk), .RN(n4306), .QN(n1254) );
  DFFRX1 \tag_r_reg[1][8]  ( .D(n3817), .CK(clk), .RN(n4306), .QN(n1255) );
  DFFRX1 \tag_r_reg[1][7]  ( .D(n3818), .CK(clk), .RN(n4306), .QN(n1256) );
  DFFRX1 \tag_r_reg[1][5]  ( .D(n3820), .CK(clk), .RN(n4306), .QN(n1258) );
  DFFRX1 \tag_r_reg[1][23]  ( .D(n3802), .CK(clk), .RN(n4307), .QN(n1240) );
  DFFRX1 \tag_r_reg[1][22]  ( .D(n3803), .CK(clk), .RN(n4307), .QN(n1241) );
  DFFRX1 \tag_r_reg[1][21]  ( .D(n3804), .CK(clk), .RN(n4307), .QN(n1242) );
  DFFRX1 \tag_r_reg[1][20]  ( .D(n3805), .CK(clk), .RN(n4307), .QN(n1243) );
  DFFRX1 \tag_r_reg[1][19]  ( .D(n3806), .CK(clk), .RN(n4307), .QN(n1244) );
  DFFRX1 \valid_r_reg[2]  ( .D(n3981), .CK(clk), .RN(n4308), .QN(n48) );
  DFFRX1 \dirty_r_reg[2]  ( .D(n3986), .CK(clk), .RN(n4309), .QN(n40) );
  DFFRX1 \valid_r_reg[0]  ( .D(n3983), .CK(clk), .RN(n4307), .QN(n50) );
  DFFRX1 \dirty_r_reg[0]  ( .D(n3984), .CK(clk), .RN(n4309), .QN(n42) );
  DFFRX1 \valid_r_reg[3]  ( .D(n3980), .CK(clk), .RN(n4308), .QN(n47) );
  DFFRX1 \dirty_r_reg[3]  ( .D(n3987), .CK(clk), .RN(n4308), .QN(n39) );
  DFFRX1 \tag_r_reg[4][23]  ( .D(n3877), .CK(clk), .RN(n4301), .QN(n1165) );
  DFFRX1 \tag_r_reg[4][22]  ( .D(n3878), .CK(clk), .RN(n4301), .QN(n1166) );
  DFFRX1 \tag_r_reg[4][21]  ( .D(n3879), .CK(clk), .RN(n4301), .QN(n1167) );
  DFFRX1 \tag_r_reg[4][20]  ( .D(n3880), .CK(clk), .RN(n4301), .QN(n1168) );
  DFFRX1 \tag_r_reg[4][19]  ( .D(n3881), .CK(clk), .RN(n4301), .QN(n1169) );
  DFFRX1 \tag_r_reg[4][11]  ( .D(n3889), .CK(clk), .RN(n4300), .QN(n1177) );
  DFFRX1 \tag_r_reg[4][10]  ( .D(n3890), .CK(clk), .RN(n4300), .QN(n1178) );
  DFFRX1 \tag_r_reg[4][9]  ( .D(n3891), .CK(clk), .RN(n4300), .QN(n1179) );
  DFFRX1 \tag_r_reg[4][8]  ( .D(n3892), .CK(clk), .RN(n4300), .QN(n1180) );
  DFFRX1 \tag_r_reg[4][7]  ( .D(n3893), .CK(clk), .RN(n4300), .QN(n1181) );
  DFFRX1 \tag_r_reg[4][5]  ( .D(n3895), .CK(clk), .RN(n4300), .QN(n1183) );
  DFFRX1 \tag_r_reg[7][23]  ( .D(n3952), .CK(clk), .RN(n4295), .QN(n1090) );
  DFFRX1 \tag_r_reg[7][22]  ( .D(n3953), .CK(clk), .RN(n4295), .QN(n1091) );
  DFFRX1 \tag_r_reg[7][21]  ( .D(n3954), .CK(clk), .RN(n4295), .QN(n1092) );
  DFFRX1 \tag_r_reg[7][20]  ( .D(n3955), .CK(clk), .RN(n4295), .QN(n1093) );
  DFFRX1 \tag_r_reg[7][19]  ( .D(n3956), .CK(clk), .RN(n4294), .QN(n1094) );
  DFFRX1 \tag_r_reg[7][16]  ( .D(n3959), .CK(clk), .RN(n4294), .QN(n1097) );
  DFFRX1 \tag_r_reg[7][10]  ( .D(n3965), .CK(clk), .RN(n4294), .QN(n1103) );
  DFFRX1 \tag_r_reg[7][9]  ( .D(n3966), .CK(clk), .RN(n4294), .QN(n1104) );
  DFFRX1 \tag_r_reg[7][8]  ( .D(n3967), .CK(clk), .RN(n4294), .QN(n1105) );
  DFFRX1 \tag_r_reg[7][7]  ( .D(n3968), .CK(clk), .RN(n4293), .QN(n1106) );
  DFFRX1 \tag_r_reg[7][5]  ( .D(n3970), .CK(clk), .RN(n4293), .QN(n1108) );
  DFFRX1 \tag_r_reg[6][23]  ( .D(n3927), .CK(clk), .RN(n4297), .QN(n1115) );
  DFFRX1 \tag_r_reg[6][22]  ( .D(n3928), .CK(clk), .RN(n4297), .QN(n1116) );
  DFFRX1 \tag_r_reg[6][21]  ( .D(n3929), .CK(clk), .RN(n4297), .QN(n1117) );
  DFFRX1 \tag_r_reg[6][20]  ( .D(n3930), .CK(clk), .RN(n4297), .QN(n1118) );
  DFFRX1 \tag_r_reg[6][19]  ( .D(n3931), .CK(clk), .RN(n4297), .QN(n1119) );
  DFFRX1 \tag_r_reg[6][11]  ( .D(n3939), .CK(clk), .RN(n4296), .QN(n1127) );
  DFFRX1 \tag_r_reg[6][10]  ( .D(n3940), .CK(clk), .RN(n4296), .QN(n1128) );
  DFFRX1 \tag_r_reg[6][9]  ( .D(n3941), .CK(clk), .RN(n4296), .QN(n1129) );
  DFFRX1 \tag_r_reg[6][8]  ( .D(n3942), .CK(clk), .RN(n4296), .QN(n1130) );
  DFFRX1 \tag_r_reg[6][7]  ( .D(n3943), .CK(clk), .RN(n4296), .QN(n1131) );
  DFFRX1 \tag_r_reg[6][5]  ( .D(n3945), .CK(clk), .RN(n4295), .QN(n1133) );
  DFFRX1 \tag_r_reg[5][23]  ( .D(n3902), .CK(clk), .RN(n4299), .QN(n1140) );
  DFFRX1 \tag_r_reg[5][22]  ( .D(n3903), .CK(clk), .RN(n4299), .QN(n1141) );
  DFFRX1 \tag_r_reg[5][21]  ( .D(n3904), .CK(clk), .RN(n4299), .QN(n1142) );
  DFFRX1 \tag_r_reg[5][20]  ( .D(n3905), .CK(clk), .RN(n4299), .QN(n1143) );
  DFFRX1 \tag_r_reg[5][19]  ( .D(n3906), .CK(clk), .RN(n4299), .QN(n1144) );
  DFFRX1 \tag_r_reg[5][11]  ( .D(n3914), .CK(clk), .RN(n4298), .QN(n1152) );
  DFFRX1 \tag_r_reg[5][10]  ( .D(n3915), .CK(clk), .RN(n4298), .QN(n1153) );
  DFFRX1 \tag_r_reg[5][9]  ( .D(n3916), .CK(clk), .RN(n4298), .QN(n1154) );
  DFFRX1 \tag_r_reg[5][8]  ( .D(n3917), .CK(clk), .RN(n4298), .QN(n1155) );
  DFFRX1 \tag_r_reg[5][7]  ( .D(n3918), .CK(clk), .RN(n4298), .QN(n1156) );
  DFFRX1 \tag_r_reg[5][5]  ( .D(n3920), .CK(clk), .RN(n4297), .QN(n1158) );
  DFFRX1 \valid_r_reg[1]  ( .D(n3982), .CK(clk), .RN(n4308), .QN(n49) );
  DFFRX1 \dirty_r_reg[1]  ( .D(n3985), .CK(clk), .RN(n4309), .QN(n41) );
  DFFRX1 \block_r_reg[1][17]  ( .D(n3631), .CK(clk), .RN(n4290), .QN(n943) );
  DFFRX1 \block_r_reg[1][16]  ( .D(n3632), .CK(clk), .RN(n4290), .QN(n944) );
  DFFRX1 \block_r_reg[1][15]  ( .D(n3633), .CK(clk), .RN(n4289), .QN(n945) );
  DFFRX1 \block_r_reg[1][14]  ( .D(n3634), .CK(clk), .RN(n4288), .QN(n946) );
  DFFRX1 \block_r_reg[1][13]  ( .D(n3635), .CK(clk), .RN(n4288), .QN(n947) );
  DFFRX1 \block_r_reg[1][12]  ( .D(n3636), .CK(clk), .RN(n4287), .QN(n948) );
  DFFRX1 \block_r_reg[1][11]  ( .D(n3637), .CK(clk), .RN(n4286), .QN(n949) );
  DFFRX1 \block_r_reg[1][10]  ( .D(n3638), .CK(clk), .RN(n4286), .QN(n950) );
  DFFRX1 \block_r_reg[4][29]  ( .D(n3235), .CK(clk), .RN(n4213), .QN(n547) );
  DFFRX1 \block_r_reg[4][28]  ( .D(n3236), .CK(clk), .RN(n4212), .QN(n548) );
  DFFRX1 \block_r_reg[4][27]  ( .D(n3237), .CK(clk), .RN(n4212), .QN(n549) );
  DFFRX1 \block_r_reg[4][26]  ( .D(n3238), .CK(clk), .RN(n4211), .QN(n550) );
  DFFRX1 \block_r_reg[4][25]  ( .D(n3239), .CK(clk), .RN(n4210), .QN(n551) );
  DFFRX1 \block_r_reg[4][24]  ( .D(n3240), .CK(clk), .RN(n4210), .QN(n552) );
  DFFRX1 \block_r_reg[4][23]  ( .D(n3241), .CK(clk), .RN(n4209), .QN(n553) );
  DFFRX1 \block_r_reg[4][22]  ( .D(n3242), .CK(clk), .RN(n4208), .QN(n554) );
  NAND2X1 U3 ( .A(n1337), .B(n4129), .Y(n1) );
  AND3X2 U4 ( .A(proc_addr[3]), .B(proc_addr[2]), .C(mem_addr[2]), .Y(n1299)
         );
  NAND2X1 U5 ( .A(n1337), .B(n1577), .Y(n2) );
  CLKBUFX2 U6 ( .A(n1699), .Y(n4057) );
  NAND2X1 U7 ( .A(n1337), .B(n1551), .Y(n3) );
  NAND2X1 U8 ( .A(n1337), .B(n1553), .Y(n4) );
  NAND2X1 U9 ( .A(n1337), .B(n1299), .Y(n5) );
  NAND2X1 U10 ( .A(n1337), .B(n1549), .Y(n6) );
  NAND2X1 U11 ( .A(n1337), .B(n4139), .Y(n7) );
  NAND2X1 U12 ( .A(n1337), .B(n4119), .Y(n8) );
  NAND2X1 U13 ( .A(proc_addr_1), .B(n4354), .Y(n9) );
  NAND2X1 U14 ( .A(proc_addr_0), .B(n4355), .Y(n10) );
  NAND2X1 U15 ( .A(n1548), .B(n1553), .Y(n11) );
  NAND2X1 U16 ( .A(n1548), .B(n1551), .Y(n12) );
  NAND2X1 U17 ( .A(n1548), .B(n1577), .Y(n13) );
  NAND2X1 U18 ( .A(n4419), .B(n64), .Y(n14) );
  OA22X1 U19 ( .A0(n4000), .A1(n1317), .B0(n2627), .B1(n14), .Y(n15) );
  NAND2X1 U20 ( .A(proc_addr_1), .B(proc_addr_0), .Y(n16) );
  OA22X1 U21 ( .A0(n4000), .A1(n1327), .B0(n2703), .B1(n4001), .Y(n17) );
  OA22X1 U22 ( .A0(n4000), .A1(n1328), .B0(n2698), .B1(n4001), .Y(n18) );
  OA22X1 U23 ( .A0(n4000), .A1(n1329), .B0(n2693), .B1(n4002), .Y(n19) );
  OA22X1 U24 ( .A0(n4000), .A1(n1330), .B0(n2688), .B1(n4002), .Y(n20) );
  OA22X1 U25 ( .A0(n4000), .A1(n1331), .B0(n2683), .B1(n4002), .Y(n21) );
  OA22X1 U26 ( .A0(n4000), .A1(n1334), .B0(n2668), .B1(n4001), .Y(n22) );
  OA22X1 U27 ( .A0(n4000), .A1(n1310), .B0(n2663), .B1(n4002), .Y(n23) );
  OA22X1 U28 ( .A0(n4000), .A1(n1332), .B0(n2678), .B1(n4002), .Y(n24) );
  OA22X1 U29 ( .A0(n4000), .A1(n1333), .B0(n2673), .B1(n4002), .Y(n25) );
  INVX12 U30 ( .A(n1524), .Y(mem_wdata[0]) );
  NOR4X2 U31 ( .A(n2623), .B(n2624), .C(n2625), .D(n2626), .Y(n1524) );
  INVX12 U32 ( .A(n1395), .Y(mem_wdata[100]) );
  NOR4X2 U33 ( .A(n2619), .B(n2620), .C(n2621), .D(n2622), .Y(n1395) );
  INVX12 U34 ( .A(n1390), .Y(mem_wdata[101]) );
  NOR4X2 U35 ( .A(n2615), .B(n2616), .C(n2617), .D(n2618), .Y(n1390) );
  INVX12 U36 ( .A(n1385), .Y(mem_wdata[102]) );
  NOR4X2 U37 ( .A(n2611), .B(n2612), .C(n2613), .D(n2614), .Y(n1385) );
  INVX12 U38 ( .A(n1380), .Y(mem_wdata[103]) );
  NOR4X2 U39 ( .A(n2607), .B(n2608), .C(n2609), .D(n2610), .Y(n1380) );
  INVX12 U40 ( .A(n1375), .Y(mem_wdata[104]) );
  NOR4X2 U41 ( .A(n2603), .B(n2604), .C(n2605), .D(n2606), .Y(n1375) );
  INVX12 U42 ( .A(n1369), .Y(mem_wdata[105]) );
  NOR4X2 U43 ( .A(n2599), .B(n2600), .C(n2601), .D(n2602), .Y(n1369) );
  INVX12 U44 ( .A(n1520), .Y(mem_wdata[106]) );
  NOR4X2 U45 ( .A(n2595), .B(n2596), .C(n2597), .D(n2598), .Y(n1520) );
  INVX12 U46 ( .A(n1515), .Y(mem_wdata[107]) );
  NOR4X2 U47 ( .A(n2591), .B(n2592), .C(n2593), .D(n2594), .Y(n1515) );
  INVX12 U48 ( .A(n1510), .Y(mem_wdata[108]) );
  NOR4X2 U49 ( .A(n2587), .B(n2588), .C(n2589), .D(n2590), .Y(n1510) );
  INVX12 U50 ( .A(n1505), .Y(mem_wdata[109]) );
  NOR4X2 U51 ( .A(n2583), .B(n2584), .C(n2585), .D(n2586), .Y(n1505) );
  INVX12 U52 ( .A(n1519), .Y(mem_wdata[10]) );
  NOR4X2 U53 ( .A(n2579), .B(n2580), .C(n2581), .D(n2582), .Y(n1519) );
  INVX12 U54 ( .A(n1500), .Y(mem_wdata[110]) );
  NOR4X2 U55 ( .A(n2575), .B(n2576), .C(n2577), .D(n2578), .Y(n1500) );
  INVX12 U56 ( .A(n1495), .Y(mem_wdata[111]) );
  NOR4X2 U57 ( .A(n2571), .B(n2572), .C(n2573), .D(n2574), .Y(n1495) );
  INVX12 U58 ( .A(n1490), .Y(mem_wdata[112]) );
  NOR4X2 U59 ( .A(n2567), .B(n2568), .C(n2569), .D(n2570), .Y(n1490) );
  INVX12 U60 ( .A(n1485), .Y(mem_wdata[113]) );
  NOR4X2 U61 ( .A(n2563), .B(n2564), .C(n2565), .D(n2566), .Y(n1485) );
  INVX12 U62 ( .A(n1480), .Y(mem_wdata[114]) );
  NOR4X2 U63 ( .A(n2559), .B(n2560), .C(n2561), .D(n2562), .Y(n1480) );
  INVX12 U64 ( .A(n1475), .Y(mem_wdata[115]) );
  NOR4X2 U65 ( .A(n2555), .B(n2556), .C(n2557), .D(n2558), .Y(n1475) );
  INVX12 U66 ( .A(n1465), .Y(mem_wdata[116]) );
  NOR4X2 U67 ( .A(n2551), .B(n2552), .C(n2553), .D(n2554), .Y(n1465) );
  INVX12 U68 ( .A(n1460), .Y(mem_wdata[117]) );
  NOR4X2 U69 ( .A(n2547), .B(n2548), .C(n2549), .D(n2550), .Y(n1460) );
  INVX12 U70 ( .A(n1455), .Y(mem_wdata[118]) );
  NOR4X2 U71 ( .A(n2543), .B(n2544), .C(n2545), .D(n2546), .Y(n1455) );
  INVX12 U72 ( .A(n1450), .Y(mem_wdata[119]) );
  NOR4X2 U73 ( .A(n2539), .B(n2540), .C(n2541), .D(n2542), .Y(n1450) );
  INVX12 U74 ( .A(n1514), .Y(mem_wdata[11]) );
  NOR4X2 U75 ( .A(n2535), .B(n2536), .C(n2537), .D(n2538), .Y(n1514) );
  INVX12 U76 ( .A(n1445), .Y(mem_wdata[120]) );
  NOR4X2 U77 ( .A(n2531), .B(n2532), .C(n2533), .D(n2534), .Y(n1445) );
  INVX12 U78 ( .A(n1440), .Y(mem_wdata[121]) );
  NOR4X2 U79 ( .A(n2527), .B(n2528), .C(n2529), .D(n2530), .Y(n1440) );
  INVX12 U80 ( .A(n1435), .Y(mem_wdata[122]) );
  NOR4X2 U81 ( .A(n2523), .B(n2524), .C(n2525), .D(n2526), .Y(n1435) );
  INVX12 U82 ( .A(n1430), .Y(mem_wdata[123]) );
  NOR4X2 U83 ( .A(n2519), .B(n2520), .C(n2521), .D(n2522), .Y(n1430) );
  INVX12 U84 ( .A(n1425), .Y(mem_wdata[124]) );
  NOR4X2 U85 ( .A(n2515), .B(n2516), .C(n2517), .D(n2518), .Y(n1425) );
  INVX12 U86 ( .A(n1420), .Y(mem_wdata[125]) );
  NOR4X2 U87 ( .A(n2511), .B(n2512), .C(n2513), .D(n2514), .Y(n1420) );
  INVX12 U88 ( .A(n1410), .Y(mem_wdata[126]) );
  NOR4X2 U89 ( .A(n2507), .B(n2508), .C(n2509), .D(n2510), .Y(n1410) );
  INVX12 U90 ( .A(n1405), .Y(mem_wdata[127]) );
  NOR4X2 U91 ( .A(n2503), .B(n2504), .C(n2505), .D(n2506), .Y(n1405) );
  INVX12 U92 ( .A(n1509), .Y(mem_wdata[12]) );
  NOR4X2 U93 ( .A(n2499), .B(n2500), .C(n2501), .D(n2502), .Y(n1509) );
  INVX12 U94 ( .A(n1504), .Y(mem_wdata[13]) );
  NOR4X2 U95 ( .A(n2495), .B(n2496), .C(n2497), .D(n2498), .Y(n1504) );
  INVX12 U96 ( .A(n1499), .Y(mem_wdata[14]) );
  NOR4X2 U97 ( .A(n2491), .B(n2492), .C(n2493), .D(n2494), .Y(n1499) );
  INVX12 U98 ( .A(n1494), .Y(mem_wdata[15]) );
  NOR4X2 U99 ( .A(n2487), .B(n2488), .C(n2489), .D(n2490), .Y(n1494) );
  INVX12 U100 ( .A(n1489), .Y(mem_wdata[16]) );
  NOR4X2 U101 ( .A(n2483), .B(n2484), .C(n2485), .D(n2486), .Y(n1489) );
  INVX12 U102 ( .A(n1484), .Y(mem_wdata[17]) );
  NOR4X2 U103 ( .A(n2479), .B(n2480), .C(n2481), .D(n2482), .Y(n1484) );
  INVX12 U104 ( .A(n1479), .Y(mem_wdata[18]) );
  NOR4X2 U105 ( .A(n2475), .B(n2476), .C(n2477), .D(n2478), .Y(n1479) );
  INVX12 U106 ( .A(n1474), .Y(mem_wdata[19]) );
  NOR4X2 U107 ( .A(n2471), .B(n2472), .C(n2473), .D(n2474), .Y(n1474) );
  INVX12 U108 ( .A(n1469), .Y(mem_wdata[1]) );
  NOR4X2 U109 ( .A(n2467), .B(n2468), .C(n2469), .D(n2470), .Y(n1469) );
  INVX12 U110 ( .A(n1464), .Y(mem_wdata[20]) );
  NOR4X2 U111 ( .A(n2463), .B(n2464), .C(n2465), .D(n2466), .Y(n1464) );
  INVX12 U112 ( .A(n1459), .Y(mem_wdata[21]) );
  NOR4X2 U113 ( .A(n2459), .B(n2460), .C(n2461), .D(n2462), .Y(n1459) );
  INVX12 U114 ( .A(n1454), .Y(mem_wdata[22]) );
  NOR4X2 U115 ( .A(n2455), .B(n2456), .C(n2457), .D(n2458), .Y(n1454) );
  INVX12 U116 ( .A(n1449), .Y(mem_wdata[23]) );
  NOR4X2 U117 ( .A(n2451), .B(n2452), .C(n2453), .D(n2454), .Y(n1449) );
  INVX12 U118 ( .A(n1444), .Y(mem_wdata[24]) );
  NOR4X2 U119 ( .A(n2447), .B(n2448), .C(n2449), .D(n2450), .Y(n1444) );
  INVX12 U120 ( .A(n1439), .Y(mem_wdata[25]) );
  NOR4X2 U121 ( .A(n2443), .B(n2444), .C(n2445), .D(n2446), .Y(n1439) );
  INVX12 U122 ( .A(n1434), .Y(mem_wdata[26]) );
  NOR4X2 U123 ( .A(n2439), .B(n2440), .C(n2441), .D(n2442), .Y(n1434) );
  INVX12 U124 ( .A(n1429), .Y(mem_wdata[27]) );
  NOR4X2 U125 ( .A(n2435), .B(n2436), .C(n2437), .D(n2438), .Y(n1429) );
  INVX12 U126 ( .A(n1424), .Y(mem_wdata[28]) );
  NOR4X2 U127 ( .A(n2431), .B(n2432), .C(n2433), .D(n2434), .Y(n1424) );
  INVX12 U128 ( .A(n1419), .Y(mem_wdata[29]) );
  NOR4X2 U129 ( .A(n2427), .B(n2428), .C(n2429), .D(n2430), .Y(n1419) );
  INVX12 U130 ( .A(n1414), .Y(mem_wdata[2]) );
  NOR4X2 U131 ( .A(n2423), .B(n2424), .C(n2425), .D(n2426), .Y(n1414) );
  INVX12 U132 ( .A(n1409), .Y(mem_wdata[30]) );
  NOR4X2 U133 ( .A(n2419), .B(n2420), .C(n2421), .D(n2422), .Y(n1409) );
  INVX12 U134 ( .A(n1404), .Y(mem_wdata[31]) );
  NOR4X2 U135 ( .A(n2415), .B(n2416), .C(n2417), .D(n2418), .Y(n1404) );
  INVX12 U136 ( .A(n1522), .Y(mem_wdata[32]) );
  NOR4X2 U137 ( .A(n2411), .B(n2412), .C(n2413), .D(n2414), .Y(n1522) );
  INVX12 U138 ( .A(n1467), .Y(mem_wdata[33]) );
  NOR4X2 U139 ( .A(n2407), .B(n2408), .C(n2409), .D(n2410), .Y(n1467) );
  INVX12 U140 ( .A(n1412), .Y(mem_wdata[34]) );
  NOR4X2 U141 ( .A(n2403), .B(n2404), .C(n2405), .D(n2406), .Y(n1412) );
  INVX12 U142 ( .A(n1397), .Y(mem_wdata[35]) );
  NOR4X2 U143 ( .A(n2399), .B(n2400), .C(n2401), .D(n2402), .Y(n1397) );
  INVX12 U144 ( .A(n1392), .Y(mem_wdata[36]) );
  NOR4X2 U145 ( .A(n2395), .B(n2396), .C(n2397), .D(n2398), .Y(n1392) );
  INVX12 U146 ( .A(n1387), .Y(mem_wdata[37]) );
  NOR4X2 U147 ( .A(n2391), .B(n2392), .C(n2393), .D(n2394), .Y(n1387) );
  INVX12 U148 ( .A(n1382), .Y(mem_wdata[38]) );
  NOR4X2 U149 ( .A(n2387), .B(n2388), .C(n2389), .D(n2390), .Y(n1382) );
  INVX12 U150 ( .A(n1377), .Y(mem_wdata[39]) );
  NOR4X2 U151 ( .A(n2383), .B(n2384), .C(n2385), .D(n2386), .Y(n1377) );
  INVX12 U152 ( .A(n1399), .Y(mem_wdata[3]) );
  NOR4X2 U153 ( .A(n2379), .B(n2380), .C(n2381), .D(n2382), .Y(n1399) );
  INVX12 U154 ( .A(n1372), .Y(mem_wdata[40]) );
  NOR4X2 U155 ( .A(n2375), .B(n2376), .C(n2377), .D(n2378), .Y(n1372) );
  INVX12 U156 ( .A(n1364), .Y(mem_wdata[41]) );
  NOR4X2 U157 ( .A(n2371), .B(n2372), .C(n2373), .D(n2374), .Y(n1364) );
  INVX12 U158 ( .A(n1517), .Y(mem_wdata[42]) );
  NOR4X2 U159 ( .A(n2367), .B(n2368), .C(n2369), .D(n2370), .Y(n1517) );
  INVX12 U160 ( .A(n1512), .Y(mem_wdata[43]) );
  NOR4X2 U161 ( .A(n2363), .B(n2364), .C(n2365), .D(n2366), .Y(n1512) );
  INVX12 U162 ( .A(n1507), .Y(mem_wdata[44]) );
  NOR4X2 U163 ( .A(n2359), .B(n2360), .C(n2361), .D(n2362), .Y(n1507) );
  INVX12 U164 ( .A(n1502), .Y(mem_wdata[45]) );
  NOR4X2 U165 ( .A(n2355), .B(n2356), .C(n2357), .D(n2358), .Y(n1502) );
  INVX12 U166 ( .A(n1497), .Y(mem_wdata[46]) );
  NOR4X2 U167 ( .A(n2351), .B(n2352), .C(n2353), .D(n2354), .Y(n1497) );
  INVX12 U168 ( .A(n1492), .Y(mem_wdata[47]) );
  NOR4X2 U169 ( .A(n2347), .B(n2348), .C(n2349), .D(n2350), .Y(n1492) );
  INVX12 U170 ( .A(n1487), .Y(mem_wdata[48]) );
  NOR4X2 U171 ( .A(n2343), .B(n2344), .C(n2345), .D(n2346), .Y(n1487) );
  INVX12 U172 ( .A(n1482), .Y(mem_wdata[49]) );
  NOR4X2 U173 ( .A(n2339), .B(n2340), .C(n2341), .D(n2342), .Y(n1482) );
  INVX12 U174 ( .A(n1394), .Y(mem_wdata[4]) );
  NOR4X2 U175 ( .A(n2335), .B(n2336), .C(n2337), .D(n2338), .Y(n1394) );
  INVX12 U176 ( .A(n1477), .Y(mem_wdata[50]) );
  NOR4X2 U177 ( .A(n2331), .B(n2332), .C(n2333), .D(n2334), .Y(n1477) );
  INVX12 U178 ( .A(n1472), .Y(mem_wdata[51]) );
  NOR4X2 U179 ( .A(n2327), .B(n2328), .C(n2329), .D(n2330), .Y(n1472) );
  INVX12 U180 ( .A(n1462), .Y(mem_wdata[52]) );
  NOR4X2 U181 ( .A(n2323), .B(n2324), .C(n2325), .D(n2326), .Y(n1462) );
  INVX12 U182 ( .A(n1457), .Y(mem_wdata[53]) );
  NOR4X2 U183 ( .A(n2319), .B(n2320), .C(n2321), .D(n2322), .Y(n1457) );
  INVX12 U184 ( .A(n1452), .Y(mem_wdata[54]) );
  NOR4X2 U185 ( .A(n2315), .B(n2316), .C(n2317), .D(n2318), .Y(n1452) );
  INVX12 U186 ( .A(n1447), .Y(mem_wdata[55]) );
  NOR4X2 U187 ( .A(n2311), .B(n2312), .C(n2313), .D(n2314), .Y(n1447) );
  INVX12 U188 ( .A(n1442), .Y(mem_wdata[56]) );
  NOR4X2 U189 ( .A(n2307), .B(n2308), .C(n2309), .D(n2310), .Y(n1442) );
  INVX12 U190 ( .A(n1437), .Y(mem_wdata[57]) );
  NOR4X2 U191 ( .A(n2303), .B(n2304), .C(n2305), .D(n2306), .Y(n1437) );
  INVX12 U192 ( .A(n1432), .Y(mem_wdata[58]) );
  NOR4X2 U193 ( .A(n2299), .B(n2300), .C(n2301), .D(n2302), .Y(n1432) );
  INVX12 U194 ( .A(n1427), .Y(mem_wdata[59]) );
  NOR4X2 U195 ( .A(n2295), .B(n2296), .C(n2297), .D(n2298), .Y(n1427) );
  INVX12 U196 ( .A(n1389), .Y(mem_wdata[5]) );
  NOR4X2 U197 ( .A(n2291), .B(n2292), .C(n2293), .D(n2294), .Y(n1389) );
  INVX12 U198 ( .A(n1422), .Y(mem_wdata[60]) );
  NOR4X2 U199 ( .A(n2287), .B(n2288), .C(n2289), .D(n2290), .Y(n1422) );
  INVX12 U200 ( .A(n1417), .Y(mem_wdata[61]) );
  NOR4X2 U201 ( .A(n2283), .B(n2284), .C(n2285), .D(n2286), .Y(n1417) );
  INVX12 U202 ( .A(n1407), .Y(mem_wdata[62]) );
  NOR4X2 U203 ( .A(n2279), .B(n2280), .C(n2281), .D(n2282), .Y(n1407) );
  INVX12 U204 ( .A(n1402), .Y(mem_wdata[63]) );
  NOR4X2 U205 ( .A(n2275), .B(n2276), .C(n2277), .D(n2278), .Y(n1402) );
  INVX12 U206 ( .A(n1521), .Y(mem_wdata[64]) );
  NOR4X2 U207 ( .A(n2271), .B(n2272), .C(n2273), .D(n2274), .Y(n1521) );
  INVX12 U208 ( .A(n1466), .Y(mem_wdata[65]) );
  NOR4X2 U209 ( .A(n2267), .B(n2268), .C(n2269), .D(n2270), .Y(n1466) );
  INVX12 U210 ( .A(n1411), .Y(mem_wdata[66]) );
  NOR4X2 U211 ( .A(n2263), .B(n2264), .C(n2265), .D(n2266), .Y(n1411) );
  INVX12 U212 ( .A(n1396), .Y(mem_wdata[67]) );
  NOR4X2 U213 ( .A(n2259), .B(n2260), .C(n2261), .D(n2262), .Y(n1396) );
  INVX12 U214 ( .A(n1391), .Y(mem_wdata[68]) );
  NOR4X2 U215 ( .A(n2255), .B(n2256), .C(n2257), .D(n2258), .Y(n1391) );
  INVX12 U216 ( .A(n1386), .Y(mem_wdata[69]) );
  NOR4X2 U217 ( .A(n2251), .B(n2252), .C(n2253), .D(n2254), .Y(n1386) );
  INVX12 U218 ( .A(n1384), .Y(mem_wdata[6]) );
  NOR4X2 U219 ( .A(n2247), .B(n2248), .C(n2249), .D(n2250), .Y(n1384) );
  INVX12 U220 ( .A(n1381), .Y(mem_wdata[70]) );
  NOR4X2 U221 ( .A(n2243), .B(n2244), .C(n2245), .D(n2246), .Y(n1381) );
  INVX12 U222 ( .A(n1376), .Y(mem_wdata[71]) );
  NOR4X2 U223 ( .A(n2239), .B(n2240), .C(n2241), .D(n2242), .Y(n1376) );
  INVX12 U224 ( .A(n1371), .Y(mem_wdata[72]) );
  NOR4X2 U225 ( .A(n2235), .B(n2236), .C(n2237), .D(n2238), .Y(n1371) );
  INVX12 U226 ( .A(n1362), .Y(mem_wdata[73]) );
  NOR4X2 U227 ( .A(n2231), .B(n2232), .C(n2233), .D(n2234), .Y(n1362) );
  INVX12 U228 ( .A(n1516), .Y(mem_wdata[74]) );
  NOR4X2 U229 ( .A(n2227), .B(n2228), .C(n2229), .D(n2230), .Y(n1516) );
  INVX12 U230 ( .A(n1511), .Y(mem_wdata[75]) );
  NOR4X2 U231 ( .A(n2223), .B(n2224), .C(n2225), .D(n2226), .Y(n1511) );
  INVX12 U232 ( .A(n1506), .Y(mem_wdata[76]) );
  NOR4X2 U233 ( .A(n2219), .B(n2220), .C(n2221), .D(n2222), .Y(n1506) );
  INVX12 U234 ( .A(n1501), .Y(mem_wdata[77]) );
  NOR4X2 U235 ( .A(n2215), .B(n2216), .C(n2217), .D(n2218), .Y(n1501) );
  INVX12 U236 ( .A(n1496), .Y(mem_wdata[78]) );
  NOR4X2 U237 ( .A(n2211), .B(n2212), .C(n2213), .D(n2214), .Y(n1496) );
  INVX12 U238 ( .A(n1491), .Y(mem_wdata[79]) );
  NOR4X2 U239 ( .A(n2207), .B(n2208), .C(n2209), .D(n2210), .Y(n1491) );
  INVX12 U240 ( .A(n1379), .Y(mem_wdata[7]) );
  NOR4X2 U241 ( .A(n2203), .B(n2204), .C(n2205), .D(n2206), .Y(n1379) );
  INVX12 U242 ( .A(n1486), .Y(mem_wdata[80]) );
  NOR4X2 U243 ( .A(n2199), .B(n2200), .C(n2201), .D(n2202), .Y(n1486) );
  INVX12 U244 ( .A(n1481), .Y(mem_wdata[81]) );
  NOR4X2 U245 ( .A(n2195), .B(n2196), .C(n2197), .D(n2198), .Y(n1481) );
  INVX12 U246 ( .A(n1476), .Y(mem_wdata[82]) );
  NOR4X2 U247 ( .A(n2191), .B(n2192), .C(n2193), .D(n2194), .Y(n1476) );
  INVX12 U248 ( .A(n1471), .Y(mem_wdata[83]) );
  NOR4X2 U249 ( .A(n2187), .B(n2188), .C(n2189), .D(n2190), .Y(n1471) );
  INVX12 U250 ( .A(n1461), .Y(mem_wdata[84]) );
  NOR4X2 U251 ( .A(n2183), .B(n2184), .C(n2185), .D(n2186), .Y(n1461) );
  INVX12 U252 ( .A(n1456), .Y(mem_wdata[85]) );
  NOR4X2 U253 ( .A(n2179), .B(n2180), .C(n2181), .D(n2182), .Y(n1456) );
  INVX12 U254 ( .A(n1451), .Y(mem_wdata[86]) );
  NOR4X2 U255 ( .A(n2175), .B(n2176), .C(n2177), .D(n2178), .Y(n1451) );
  INVX12 U256 ( .A(n1446), .Y(mem_wdata[87]) );
  NOR4X2 U257 ( .A(n2171), .B(n2172), .C(n2173), .D(n2174), .Y(n1446) );
  INVX12 U258 ( .A(n1441), .Y(mem_wdata[88]) );
  NOR4X2 U259 ( .A(n2167), .B(n2168), .C(n2169), .D(n2170), .Y(n1441) );
  INVX12 U260 ( .A(n1436), .Y(mem_wdata[89]) );
  NOR4X2 U261 ( .A(n2163), .B(n2164), .C(n2165), .D(n2166), .Y(n1436) );
  INVX12 U262 ( .A(n1374), .Y(mem_wdata[8]) );
  NOR4X2 U263 ( .A(n2159), .B(n2160), .C(n2161), .D(n2162), .Y(n1374) );
  INVX12 U264 ( .A(n1431), .Y(mem_wdata[90]) );
  NOR4X2 U265 ( .A(n2155), .B(n2156), .C(n2157), .D(n2158), .Y(n1431) );
  INVX12 U266 ( .A(n1426), .Y(mem_wdata[91]) );
  NOR4X2 U267 ( .A(n2151), .B(n2152), .C(n2153), .D(n2154), .Y(n1426) );
  INVX12 U268 ( .A(n1421), .Y(mem_wdata[92]) );
  NOR4X2 U269 ( .A(n2147), .B(n2148), .C(n2149), .D(n2150), .Y(n1421) );
  INVX12 U270 ( .A(n1416), .Y(mem_wdata[93]) );
  NOR4X2 U271 ( .A(n2143), .B(n2144), .C(n2145), .D(n2146), .Y(n1416) );
  INVX12 U272 ( .A(n1406), .Y(mem_wdata[94]) );
  NOR4X2 U273 ( .A(n2139), .B(n2140), .C(n2141), .D(n2142), .Y(n1406) );
  INVX12 U274 ( .A(n1401), .Y(mem_wdata[95]) );
  NOR4X2 U275 ( .A(n2135), .B(n2136), .C(n2137), .D(n2138), .Y(n1401) );
  INVX12 U276 ( .A(n1525), .Y(mem_wdata[96]) );
  NOR4X2 U277 ( .A(n2131), .B(n2132), .C(n2133), .D(n2134), .Y(n1525) );
  INVX12 U278 ( .A(n1470), .Y(mem_wdata[97]) );
  NOR4X2 U279 ( .A(n2127), .B(n2128), .C(n2129), .D(n2130), .Y(n1470) );
  INVX12 U280 ( .A(n1415), .Y(mem_wdata[98]) );
  NOR4X2 U281 ( .A(n2123), .B(n2124), .C(n2125), .D(n2126), .Y(n1415) );
  INVX12 U282 ( .A(n1400), .Y(mem_wdata[99]) );
  NOR4X2 U283 ( .A(n2119), .B(n2120), .C(n2121), .D(n2122), .Y(n1400) );
  INVX12 U284 ( .A(n1367), .Y(mem_wdata[9]) );
  NOR4X2 U285 ( .A(n2115), .B(n2116), .C(n2117), .D(n2118), .Y(n1367) );
  INVX12 U286 ( .A(n17), .Y(mem_addr[19]) );
  INVX12 U287 ( .A(n18), .Y(mem_addr[20]) );
  INVX12 U288 ( .A(n19), .Y(mem_addr[21]) );
  INVX12 U289 ( .A(n20), .Y(mem_addr[22]) );
  INVX12 U290 ( .A(n21), .Y(mem_addr[23]) );
  INVX12 U291 ( .A(n24), .Y(mem_addr[24]) );
  INVX12 U292 ( .A(n25), .Y(mem_addr[25]) );
  INVX12 U293 ( .A(n22), .Y(mem_addr[26]) );
  INVX12 U294 ( .A(n23), .Y(mem_addr[27]) );
  INVX12 U295 ( .A(n15), .Y(mem_addr[9]) );
  OA22X1 U296 ( .A0(n4000), .A1(n1326), .B0(n2708), .B1(n4001), .Y(n4420) );
  INVX12 U297 ( .A(n4420), .Y(mem_addr[18]) );
  OA22X1 U298 ( .A0(n4000), .A1(n1325), .B0(n2713), .B1(n4001), .Y(n4421) );
  INVX12 U299 ( .A(n4421), .Y(mem_addr[17]) );
  OA22X1 U300 ( .A0(n4000), .A1(n1324), .B0(n2718), .B1(n4001), .Y(n4422) );
  INVX12 U301 ( .A(n4422), .Y(mem_addr[16]) );
  OA22X1 U302 ( .A0(n4000), .A1(n1323), .B0(n2723), .B1(n4002), .Y(n4423) );
  INVX12 U303 ( .A(n4423), .Y(mem_addr[15]) );
  OA22X1 U304 ( .A0(n4000), .A1(n1316), .B0(n2633), .B1(n14), .Y(n4429) );
  INVX12 U305 ( .A(n4429), .Y(mem_addr[8]) );
  OA22X1 U306 ( .A0(n4000), .A1(n1322), .B0(n2728), .B1(n14), .Y(n4424) );
  INVX12 U307 ( .A(n4424), .Y(mem_addr[14]) );
  OA22X1 U308 ( .A0(n4000), .A1(n1315), .B0(n2638), .B1(n4002), .Y(n4430) );
  INVX12 U309 ( .A(n4430), .Y(mem_addr[7]) );
  OA22X1 U310 ( .A0(n4000), .A1(n1321), .B0(n2733), .B1(n4001), .Y(n4425) );
  INVX12 U311 ( .A(n4425), .Y(mem_addr[13]) );
  OA22X1 U312 ( .A0(n4000), .A1(n1313), .B0(n2648), .B1(n4001), .Y(n4432) );
  INVX12 U313 ( .A(n4432), .Y(mem_addr[5]) );
  CLKINVX1 U314 ( .A(proc_addr[4]), .Y(n1335) );
  OA22X1 U315 ( .A0(n4000), .A1(n1319), .B0(n2743), .B1(n4001), .Y(n4427) );
  INVX12 U316 ( .A(n4427), .Y(mem_addr[11]) );
  OA22X1 U317 ( .A0(n4000), .A1(n1314), .B0(n2643), .B1(n4001), .Y(n4431) );
  INVX12 U318 ( .A(n4431), .Y(mem_addr[6]) );
  OA22X1 U319 ( .A0(n4000), .A1(n1320), .B0(n2738), .B1(n4002), .Y(n4426) );
  INVX12 U320 ( .A(n4426), .Y(mem_addr[12]) );
  OA22X1 U321 ( .A0(n4000), .A1(n1312), .B0(n2653), .B1(n4002), .Y(n4433) );
  INVX12 U322 ( .A(n4433), .Y(mem_addr[4]) );
  INVX12 U323 ( .A(n1361), .Y(mem_read) );
  OA22X1 U324 ( .A0(n4000), .A1(n1318), .B0(n2748), .B1(n4002), .Y(n4428) );
  INVX12 U325 ( .A(n4428), .Y(mem_addr[10]) );
  OA22X1 U326 ( .A0(n4000), .A1(n1311), .B0(n2658), .B1(n4002), .Y(n4434) );
  INVX12 U327 ( .A(n4434), .Y(mem_addr[3]) );
  BUFX12 U328 ( .A(n4419), .Y(mem_write) );
  CLKINVX1 U329 ( .A(n4205), .Y(n4346) );
  NAND3X1 U330 ( .A(n1570), .B(n4129), .C(n1337), .Y(n1294) );
  NOR2X2 U331 ( .A(n4418), .B(n1361), .Y(n1548) );
  NOR3X1 U332 ( .A(proc_addr[3]), .B(mem_addr[2]), .C(n4358), .Y(n1549) );
  NOR3X1 U333 ( .A(proc_addr[3]), .B(mem_addr[2]), .C(proc_addr[2]), .Y(n1577)
         );
  NOR3X1 U334 ( .A(proc_addr[2]), .B(mem_addr[2]), .C(n4361), .Y(n1551) );
  OAI21XL U335 ( .A0(proc_write), .A1(n4353), .B0(n1576), .Y(n1568) );
  OAI22XL U336 ( .A0(n1552), .A1(n1238), .B0(n1550), .B1(n1213), .Y(n2661) );
  OAI22XL U337 ( .A0(n1552), .A1(n1237), .B0(n1550), .B1(n1212), .Y(n2656) );
  OAI22XL U338 ( .A0(n1558), .A1(n1236), .B0(n1550), .B1(n1211), .Y(n2651) );
  OAI22XL U339 ( .A0(n1552), .A1(n1235), .B0(n1550), .B1(n1210), .Y(n2646) );
  OAI22XL U340 ( .A0(n1552), .A1(n1226), .B0(n1550), .B1(n1201), .Y(n2726) );
  OAI22XL U341 ( .A0(n1552), .A1(n1225), .B0(n1550), .B1(n1200), .Y(n2721) );
  OAI22XL U342 ( .A0(n1558), .A1(n1224), .B0(n1550), .B1(n1199), .Y(n2716) );
  OAI22XL U343 ( .A0(n1558), .A1(n1223), .B0(n1550), .B1(n1198), .Y(n2711) );
  OAI22XL U344 ( .A0(n1558), .A1(n1222), .B0(n1550), .B1(n1197), .Y(n2706) );
  OAI22XL U345 ( .A0(n1558), .A1(n1221), .B0(n1550), .B1(n1196), .Y(n2701) );
  OAI22XL U346 ( .A0(n1558), .A1(n1220), .B0(n1550), .B1(n1195), .Y(n2696) );
  OAI22XL U347 ( .A0(n1552), .A1(n1219), .B0(n1550), .B1(n1194), .Y(n2691) );
  OAI22XL U348 ( .A0(n1552), .A1(n1218), .B0(n1550), .B1(n1193), .Y(n2686) );
  OAI22XL U349 ( .A0(n1552), .A1(n1217), .B0(n1550), .B1(n1192), .Y(n2681) );
  OAI22XL U350 ( .A0(n1552), .A1(n1216), .B0(n1550), .B1(n1191), .Y(n2676) );
  OAI22XL U351 ( .A0(n1552), .A1(n1215), .B0(n1550), .B1(n1190), .Y(n2671) );
  OAI22XL U352 ( .A0(n1558), .A1(n1214), .B0(n1550), .B1(n1189), .Y(n2666) );
  OAI22XL U353 ( .A0(n3999), .A1(n1288), .B0(n1351), .B1(n1263), .Y(n2662) );
  OAI22XL U354 ( .A0(n3999), .A1(n1287), .B0(n1355), .B1(n1262), .Y(n2657) );
  OAI22XL U355 ( .A0(n3999), .A1(n1286), .B0(n1354), .B1(n1261), .Y(n2652) );
  OAI22XL U356 ( .A0(n3999), .A1(n1285), .B0(n1350), .B1(n1260), .Y(n2647) );
  OAI22XL U357 ( .A0(n3998), .A1(n1284), .B0(n1357), .B1(n1259), .Y(n2642) );
  OAI22XL U358 ( .A0(n3998), .A1(n1283), .B0(n1357), .B1(n1258), .Y(n2637) );
  OAI22XL U359 ( .A0(n3998), .A1(n1282), .B0(n1357), .B1(n1257), .Y(n2632) );
  OAI22XL U360 ( .A0(n3999), .A1(n1276), .B0(n1355), .B1(n1251), .Y(n2727) );
  OAI22XL U361 ( .A0(n3999), .A1(n1275), .B0(n1352), .B1(n1250), .Y(n2722) );
  OAI22XL U362 ( .A0(n3999), .A1(n1274), .B0(n1351), .B1(n1249), .Y(n2717) );
  OAI22XL U363 ( .A0(n3999), .A1(n1273), .B0(n1351), .B1(n1248), .Y(n2712) );
  OAI22XL U364 ( .A0(n3999), .A1(n1272), .B0(n1351), .B1(n1247), .Y(n2707) );
  OAI22XL U365 ( .A0(n3999), .A1(n1271), .B0(n1351), .B1(n1246), .Y(n2702) );
  OAI22XL U366 ( .A0(n3999), .A1(n1270), .B0(n1354), .B1(n1245), .Y(n2697) );
  OAI22XL U367 ( .A0(n3999), .A1(n1269), .B0(n1351), .B1(n1244), .Y(n2692) );
  OAI22XL U368 ( .A0(n3999), .A1(n1268), .B0(n1351), .B1(n1243), .Y(n2687) );
  OAI22XL U369 ( .A0(n3999), .A1(n1267), .B0(n1354), .B1(n1242), .Y(n2682) );
  OAI22XL U370 ( .A0(n3999), .A1(n1266), .B0(n1351), .B1(n1241), .Y(n2677) );
  OAI22XL U371 ( .A0(n3999), .A1(n1265), .B0(n1351), .B1(n1240), .Y(n2672) );
  OAI22XL U372 ( .A0(n3999), .A1(n1264), .B0(n1351), .B1(n1239), .Y(n2667) );
  OAI22XL U373 ( .A0(n2628), .A1(n1281), .B0(n1353), .B1(n1256), .Y(n2752) );
  OAI22XL U374 ( .A0(n1701), .A1(n1234), .B0(n1546), .B1(n1209), .Y(n2641) );
  OAI22XL U375 ( .A0(n1701), .A1(n1233), .B0(n1546), .B1(n1208), .Y(n2636) );
  OAI22XL U376 ( .A0(n1701), .A1(n1232), .B0(n1546), .B1(n1207), .Y(n2631) );
  OAI22XL U377 ( .A0(n1580), .A1(n1231), .B0(n1363), .B1(n1206), .Y(n2751) );
  OAI22XL U378 ( .A0(n3998), .A1(n1088), .B0(n1357), .B1(n960), .Y(n2624) );
  OAI22XL U379 ( .A0(n1703), .A1(n1087), .B0(n1355), .B1(n959), .Y(n2468) );
  OAI22XL U380 ( .A0(n3996), .A1(n1086), .B0(n1350), .B1(n958), .Y(n2424) );
  OAI22XL U381 ( .A0(n3996), .A1(n1085), .B0(n1350), .B1(n957), .Y(n2380) );
  OAI22XL U382 ( .A0(n3998), .A1(n988), .B0(n1357), .B1(n860), .Y(n2620) );
  OAI22XL U383 ( .A0(n3995), .A1(n1084), .B0(n1357), .B1(n956), .Y(n2336) );
  OAI22XL U384 ( .A0(n3998), .A1(n987), .B0(n1357), .B1(n859), .Y(n2616) );
  OAI22XL U385 ( .A0(n3997), .A1(n1083), .B0(n1352), .B1(n955), .Y(n2292) );
  OAI22XL U386 ( .A0(n3998), .A1(n986), .B0(n1357), .B1(n858), .Y(n2612) );
  OAI22XL U387 ( .A0(n3996), .A1(n1082), .B0(n1350), .B1(n954), .Y(n2248) );
  OAI22XL U388 ( .A0(n3998), .A1(n985), .B0(n1357), .B1(n857), .Y(n2608) );
  OAI22XL U389 ( .A0(n1704), .A1(n1081), .B0(n1354), .B1(n953), .Y(n2204) );
  OAI22XL U390 ( .A0(n3998), .A1(n984), .B0(n1357), .B1(n856), .Y(n2604) );
  OAI22XL U391 ( .A0(n1704), .A1(n1080), .B0(n1354), .B1(n952), .Y(n2160) );
  OAI22XL U392 ( .A0(n3998), .A1(n983), .B0(n1357), .B1(n855), .Y(n2600) );
  OAI22XL U393 ( .A0(n3998), .A1(n982), .B0(n1357), .B1(n854), .Y(n2596) );
  OAI22XL U394 ( .A0(n3998), .A1(n1078), .B0(n1357), .B1(n950), .Y(n2580) );
  OAI22XL U395 ( .A0(n3998), .A1(n981), .B0(n1357), .B1(n853), .Y(n2592) );
  OAI22XL U396 ( .A0(n3997), .A1(n1077), .B0(n1356), .B1(n949), .Y(n2536) );
  OAI22XL U397 ( .A0(n3998), .A1(n980), .B0(n1357), .B1(n852), .Y(n2588) );
  OAI22XL U398 ( .A0(n1703), .A1(n1076), .B0(n1355), .B1(n948), .Y(n2500) );
  OAI22XL U399 ( .A0(n3998), .A1(n979), .B0(n1357), .B1(n851), .Y(n2584) );
  OAI22XL U400 ( .A0(n1703), .A1(n1075), .B0(n1355), .B1(n947), .Y(n2496) );
  OAI22XL U401 ( .A0(n3998), .A1(n978), .B0(n1357), .B1(n850), .Y(n2576) );
  OAI22XL U402 ( .A0(n1703), .A1(n1074), .B0(n1355), .B1(n946), .Y(n2492) );
  OAI22XL U403 ( .A0(n3998), .A1(n977), .B0(n1357), .B1(n849), .Y(n2572) );
  OAI22XL U404 ( .A0(n1703), .A1(n1073), .B0(n1355), .B1(n945), .Y(n2488) );
  OAI22XL U405 ( .A0(n3997), .A1(n976), .B0(n1356), .B1(n848), .Y(n2568) );
  OAI22XL U406 ( .A0(n1703), .A1(n1072), .B0(n1355), .B1(n944), .Y(n2484) );
  OAI22XL U407 ( .A0(n3997), .A1(n975), .B0(n1356), .B1(n847), .Y(n2564) );
  OAI22XL U408 ( .A0(n1703), .A1(n1071), .B0(n1355), .B1(n943), .Y(n2480) );
  OAI22XL U409 ( .A0(n3997), .A1(n974), .B0(n1356), .B1(n846), .Y(n2560) );
  OAI22XL U410 ( .A0(n1704), .A1(n1070), .B0(n1355), .B1(n942), .Y(n2476) );
  OAI22XL U411 ( .A0(n3997), .A1(n973), .B0(n1356), .B1(n845), .Y(n2556) );
  OAI22XL U412 ( .A0(n1704), .A1(n1069), .B0(n1355), .B1(n941), .Y(n2472) );
  OAI22XL U413 ( .A0(n3997), .A1(n972), .B0(n1356), .B1(n844), .Y(n2552) );
  OAI22XL U414 ( .A0(n1704), .A1(n1068), .B0(n1355), .B1(n940), .Y(n2464) );
  OAI22XL U415 ( .A0(n3997), .A1(n971), .B0(n1356), .B1(n843), .Y(n2548) );
  OAI22XL U416 ( .A0(n2628), .A1(n1067), .B0(n1355), .B1(n939), .Y(n2460) );
  OAI22XL U417 ( .A0(n3997), .A1(n970), .B0(n1356), .B1(n842), .Y(n2544) );
  OAI22XL U418 ( .A0(n1703), .A1(n1066), .B0(n1355), .B1(n938), .Y(n2456) );
  OAI22XL U419 ( .A0(n3997), .A1(n969), .B0(n1356), .B1(n841), .Y(n2540) );
  OAI22XL U420 ( .A0(n1703), .A1(n1065), .B0(n1355), .B1(n937), .Y(n2452) );
  OAI22XL U421 ( .A0(n3997), .A1(n968), .B0(n1356), .B1(n840), .Y(n2532) );
  OAI22XL U422 ( .A0(n1703), .A1(n1064), .B0(n1355), .B1(n936), .Y(n2448) );
  OAI22XL U423 ( .A0(n3997), .A1(n967), .B0(n1356), .B1(n839), .Y(n2528) );
  OAI22XL U424 ( .A0(n1703), .A1(n1063), .B0(n1355), .B1(n935), .Y(n2444) );
  OAI22XL U425 ( .A0(n3997), .A1(n966), .B0(n1356), .B1(n838), .Y(n2524) );
  OAI22XL U426 ( .A0(n1704), .A1(n1062), .B0(n1355), .B1(n934), .Y(n2440) );
  OAI22XL U427 ( .A0(n3997), .A1(n965), .B0(n1356), .B1(n837), .Y(n2520) );
  OAI22XL U428 ( .A0(n1704), .A1(n1061), .B0(n1355), .B1(n933), .Y(n2436) );
  OAI22XL U429 ( .A0(n3997), .A1(n964), .B0(n1356), .B1(n836), .Y(n2516) );
  OAI22XL U430 ( .A0(n3996), .A1(n1060), .B0(n1350), .B1(n932), .Y(n2432) );
  OAI22XL U431 ( .A0(n3997), .A1(n963), .B0(n1356), .B1(n835), .Y(n2512) );
  OAI22XL U432 ( .A0(n3996), .A1(n1059), .B0(n1350), .B1(n931), .Y(n2428) );
  OAI22XL U433 ( .A0(n3997), .A1(n962), .B0(n1356), .B1(n834), .Y(n2508) );
  OAI22XL U434 ( .A0(n3996), .A1(n1058), .B0(n1350), .B1(n930), .Y(n2420) );
  OAI22XL U435 ( .A0(n3997), .A1(n961), .B0(n1356), .B1(n833), .Y(n2504) );
  OAI22XL U436 ( .A0(n3996), .A1(n1057), .B0(n1350), .B1(n929), .Y(n2416) );
  OAI22XL U437 ( .A0(n3996), .A1(n1056), .B0(n1352), .B1(n928), .Y(n2412) );
  OAI22XL U438 ( .A0(n1704), .A1(n1024), .B0(n1351), .B1(n896), .Y(n2272) );
  OAI22XL U439 ( .A0(n3996), .A1(n1055), .B0(n1350), .B1(n927), .Y(n2408) );
  OAI22XL U440 ( .A0(n1704), .A1(n1023), .B0(n1353), .B1(n895), .Y(n2268) );
  OAI22XL U441 ( .A0(n3996), .A1(n1054), .B0(n1350), .B1(n926), .Y(n2404) );
  OAI22XL U442 ( .A0(n1703), .A1(n1022), .B0(n1350), .B1(n894), .Y(n2264) );
  OAI22XL U443 ( .A0(n3996), .A1(n1053), .B0(n1352), .B1(n925), .Y(n2400) );
  OAI22XL U444 ( .A0(n1703), .A1(n1021), .B0(n1352), .B1(n893), .Y(n2260) );
  OAI22XL U445 ( .A0(n3996), .A1(n1052), .B0(n1352), .B1(n924), .Y(n2396) );
  OAI22XL U446 ( .A0(n3995), .A1(n1020), .B0(n1352), .B1(n892), .Y(n2256) );
  OAI22XL U447 ( .A0(n3996), .A1(n1051), .B0(n1352), .B1(n923), .Y(n2392) );
  OAI22XL U448 ( .A0(n3998), .A1(n1019), .B0(n1352), .B1(n891), .Y(n2252) );
  OAI22XL U449 ( .A0(n3996), .A1(n1050), .B0(n1352), .B1(n922), .Y(n2388) );
  OAI22XL U450 ( .A0(n3998), .A1(n1018), .B0(n4356), .B1(n890), .Y(n2244) );
  OAI22XL U451 ( .A0(n3996), .A1(n1049), .B0(n1352), .B1(n921), .Y(n2384) );
  OAI22XL U452 ( .A0(n3996), .A1(n1017), .B0(n4356), .B1(n889), .Y(n2240) );
  OAI22XL U453 ( .A0(n3996), .A1(n1048), .B0(n1352), .B1(n920), .Y(n2376) );
  OAI22XL U454 ( .A0(n3997), .A1(n1016), .B0(n4356), .B1(n888), .Y(n2236) );
  OAI22XL U455 ( .A0(n3996), .A1(n1047), .B0(n1352), .B1(n919), .Y(n2372) );
  OAI22XL U456 ( .A0(n3998), .A1(n1015), .B0(n4356), .B1(n887), .Y(n2232) );
  OAI22XL U457 ( .A0(n3995), .A1(n1046), .B0(n1351), .B1(n918), .Y(n2368) );
  OAI22XL U458 ( .A0(n4360), .A1(n1014), .B0(n1354), .B1(n886), .Y(n2228) );
  OAI22XL U459 ( .A0(n3995), .A1(n1045), .B0(n1351), .B1(n917), .Y(n2364) );
  OAI22XL U460 ( .A0(n4360), .A1(n1013), .B0(n1354), .B1(n885), .Y(n2224) );
  OAI22XL U461 ( .A0(n3995), .A1(n1044), .B0(n1356), .B1(n916), .Y(n2360) );
  OAI22XL U462 ( .A0(n1704), .A1(n1012), .B0(n1354), .B1(n884), .Y(n2220) );
  OAI22XL U463 ( .A0(n3995), .A1(n1043), .B0(n1350), .B1(n915), .Y(n2356) );
  OAI22XL U464 ( .A0(n1704), .A1(n1011), .B0(n1354), .B1(n883), .Y(n2216) );
  OAI22XL U465 ( .A0(n3995), .A1(n1042), .B0(n1355), .B1(n914), .Y(n2352) );
  OAI22XL U466 ( .A0(n1704), .A1(n1010), .B0(n1354), .B1(n882), .Y(n2212) );
  OAI22XL U467 ( .A0(n3995), .A1(n1041), .B0(n1356), .B1(n913), .Y(n2348) );
  OAI22XL U468 ( .A0(n1704), .A1(n1009), .B0(n1354), .B1(n881), .Y(n2208) );
  OAI22XL U469 ( .A0(n3995), .A1(n1040), .B0(n4356), .B1(n912), .Y(n2344) );
  OAI22XL U470 ( .A0(n1704), .A1(n1008), .B0(n1354), .B1(n880), .Y(n2200) );
  OAI22XL U471 ( .A0(n3995), .A1(n1039), .B0(n1351), .B1(n911), .Y(n2340) );
  OAI22XL U472 ( .A0(n4360), .A1(n1007), .B0(n1354), .B1(n879), .Y(n2196) );
  OAI22XL U473 ( .A0(n3995), .A1(n1038), .B0(n1351), .B1(n910), .Y(n2332) );
  OAI22XL U474 ( .A0(n4360), .A1(n1006), .B0(n1354), .B1(n878), .Y(n2192) );
  OAI22XL U475 ( .A0(n3995), .A1(n1037), .B0(n1356), .B1(n909), .Y(n2328) );
  OAI22XL U476 ( .A0(n4360), .A1(n1005), .B0(n1354), .B1(n877), .Y(n2188) );
  OAI22XL U477 ( .A0(n3995), .A1(n1036), .B0(n1357), .B1(n908), .Y(n2324) );
  OAI22XL U478 ( .A0(n1704), .A1(n1004), .B0(n1354), .B1(n876), .Y(n2184) );
  OAI22XL U479 ( .A0(n3995), .A1(n1035), .B0(n1351), .B1(n907), .Y(n2320) );
  OAI22XL U480 ( .A0(n4360), .A1(n1003), .B0(n1354), .B1(n875), .Y(n2180) );
  OAI22XL U481 ( .A0(n3995), .A1(n1034), .B0(n1355), .B1(n906), .Y(n2316) );
  OAI22XL U482 ( .A0(n1704), .A1(n1002), .B0(n1354), .B1(n874), .Y(n2176) );
  OAI22XL U483 ( .A0(n3995), .A1(n1033), .B0(n1352), .B1(n905), .Y(n2312) );
  OAI22XL U484 ( .A0(n1704), .A1(n1001), .B0(n1354), .B1(n873), .Y(n2172) );
  OAI22XL U485 ( .A0(n3995), .A1(n1032), .B0(n1357), .B1(n904), .Y(n2308) );
  OAI22XL U486 ( .A0(n1704), .A1(n1000), .B0(n1354), .B1(n872), .Y(n2168) );
  OAI22XL U487 ( .A0(n3995), .A1(n1031), .B0(n1350), .B1(n903), .Y(n2304) );
  OAI22XL U488 ( .A0(n3995), .A1(n1030), .B0(n1352), .B1(n902), .Y(n2300) );
  OAI22XL U489 ( .A0(n3996), .A1(n1029), .B0(n1352), .B1(n901), .Y(n2296) );
  OAI22XL U490 ( .A0(n3995), .A1(n1028), .B0(n1352), .B1(n900), .Y(n2288) );
  OAI22XL U491 ( .A0(n3996), .A1(n1027), .B0(n1352), .B1(n899), .Y(n2284) );
  OAI22XL U492 ( .A0(n3995), .A1(n1026), .B0(n1352), .B1(n898), .Y(n2280) );
  OAI22XL U493 ( .A0(n3996), .A1(n1025), .B0(n1352), .B1(n897), .Y(n2276) );
  OAI22XL U494 ( .A0(n2628), .A1(n992), .B0(n1353), .B1(n864), .Y(n2132) );
  OAI22XL U495 ( .A0(n2628), .A1(n991), .B0(n1353), .B1(n863), .Y(n2128) );
  OAI22XL U496 ( .A0(n2628), .A1(n990), .B0(n1353), .B1(n862), .Y(n2124) );
  OAI22XL U497 ( .A0(n2628), .A1(n989), .B0(n1353), .B1(n861), .Y(n2120) );
  OAI22XL U498 ( .A0(n2628), .A1(n1079), .B0(n1353), .B1(n951), .Y(n2116) );
  OAI22XL U499 ( .A0(n2628), .A1(n999), .B0(n1353), .B1(n871), .Y(n2164) );
  OAI22XL U500 ( .A0(n2628), .A1(n998), .B0(n1353), .B1(n870), .Y(n2156) );
  OAI22XL U501 ( .A0(n2628), .A1(n997), .B0(n1353), .B1(n869), .Y(n2152) );
  OAI22XL U502 ( .A0(n2628), .A1(n996), .B0(n1353), .B1(n868), .Y(n2148) );
  OAI22XL U503 ( .A0(n2628), .A1(n995), .B0(n1353), .B1(n867), .Y(n2144) );
  OAI22XL U504 ( .A0(n2628), .A1(n994), .B0(n1353), .B1(n866), .Y(n2140) );
  OAI22XL U505 ( .A0(n2628), .A1(n993), .B0(n1353), .B1(n865), .Y(n2136) );
  OAI22XL U506 ( .A0(n2628), .A1(n42), .B0(n1353), .B1(n41), .Y(n1572) );
  OAI22XL U507 ( .A0(n4118), .A1(n1182), .B0(n4127), .B1(n1157), .Y(n2630) );
  OAI22XL U508 ( .A0(n1558), .A1(n1230), .B0(n1528), .B1(n1205), .Y(n2746) );
  OAI22XL U509 ( .A0(n1580), .A1(n1229), .B0(n1365), .B1(n1204), .Y(n2741) );
  OAI22XL U510 ( .A0(n1558), .A1(n1228), .B0(n1365), .B1(n1203), .Y(n2736) );
  OAI22XL U511 ( .A0(n1693), .A1(n1227), .B0(n1528), .B1(n1202), .Y(n2731) );
  OAI22XL U512 ( .A0(n3999), .A1(n1280), .B0(n1356), .B1(n1255), .Y(n2747) );
  OAI22XL U513 ( .A0(n3999), .A1(n1279), .B0(n1357), .B1(n1254), .Y(n2742) );
  OAI22XL U514 ( .A0(n3999), .A1(n1278), .B0(n1351), .B1(n1253), .Y(n2737) );
  OAI22XL U515 ( .A0(n3997), .A1(n1277), .B0(n1351), .B1(n1252), .Y(n2732) );
  CLKBUFX3 U516 ( .A(n4333), .Y(n4214) );
  CLKBUFX3 U517 ( .A(n4333), .Y(n4215) );
  CLKBUFX3 U518 ( .A(n4333), .Y(n4216) );
  CLKBUFX3 U519 ( .A(n4333), .Y(n4217) );
  CLKBUFX3 U520 ( .A(n4332), .Y(n4218) );
  CLKBUFX3 U521 ( .A(n4332), .Y(n4219) );
  CLKBUFX3 U522 ( .A(n4332), .Y(n4220) );
  CLKBUFX3 U523 ( .A(n4332), .Y(n4221) );
  CLKBUFX3 U524 ( .A(n4331), .Y(n4222) );
  CLKBUFX3 U525 ( .A(n4331), .Y(n4223) );
  CLKBUFX3 U526 ( .A(n4331), .Y(n4224) );
  CLKBUFX3 U527 ( .A(n4331), .Y(n4225) );
  CLKBUFX3 U528 ( .A(n4330), .Y(n4226) );
  CLKBUFX3 U529 ( .A(n4330), .Y(n4227) );
  CLKBUFX3 U530 ( .A(n4330), .Y(n4228) );
  CLKBUFX3 U531 ( .A(n4330), .Y(n4229) );
  CLKBUFX3 U532 ( .A(n4329), .Y(n4230) );
  CLKBUFX3 U533 ( .A(n4329), .Y(n4231) );
  CLKBUFX3 U534 ( .A(n4329), .Y(n4232) );
  CLKBUFX3 U535 ( .A(n4329), .Y(n4233) );
  CLKBUFX3 U536 ( .A(n4328), .Y(n4234) );
  CLKBUFX3 U537 ( .A(n4328), .Y(n4235) );
  CLKBUFX3 U538 ( .A(n4328), .Y(n4236) );
  CLKBUFX3 U539 ( .A(n4328), .Y(n4237) );
  CLKBUFX3 U540 ( .A(n4327), .Y(n4238) );
  CLKBUFX3 U541 ( .A(n4327), .Y(n4239) );
  CLKBUFX3 U542 ( .A(n4327), .Y(n4240) );
  CLKBUFX3 U543 ( .A(n4327), .Y(n4241) );
  CLKBUFX3 U544 ( .A(n4326), .Y(n4242) );
  CLKBUFX3 U545 ( .A(n4326), .Y(n4243) );
  CLKBUFX3 U546 ( .A(n4326), .Y(n4244) );
  CLKBUFX3 U547 ( .A(n4326), .Y(n4245) );
  CLKBUFX3 U548 ( .A(n4325), .Y(n4246) );
  CLKBUFX3 U549 ( .A(n4325), .Y(n4247) );
  CLKBUFX3 U550 ( .A(n4325), .Y(n4248) );
  CLKBUFX3 U551 ( .A(n4325), .Y(n4249) );
  CLKBUFX3 U552 ( .A(n4324), .Y(n4250) );
  CLKBUFX3 U553 ( .A(n4324), .Y(n4251) );
  CLKBUFX3 U554 ( .A(n4324), .Y(n4252) );
  CLKBUFX3 U555 ( .A(n4324), .Y(n4253) );
  CLKBUFX3 U556 ( .A(n4323), .Y(n4254) );
  CLKBUFX3 U557 ( .A(n4323), .Y(n4255) );
  CLKBUFX3 U558 ( .A(n4323), .Y(n4256) );
  CLKBUFX3 U559 ( .A(n4323), .Y(n4257) );
  CLKBUFX3 U560 ( .A(n4322), .Y(n4258) );
  CLKBUFX3 U561 ( .A(n4322), .Y(n4259) );
  CLKBUFX3 U562 ( .A(n4322), .Y(n4260) );
  CLKBUFX3 U563 ( .A(n4322), .Y(n4261) );
  CLKBUFX3 U564 ( .A(n4321), .Y(n4262) );
  CLKBUFX3 U565 ( .A(n4321), .Y(n4263) );
  CLKBUFX3 U566 ( .A(n4321), .Y(n4264) );
  CLKBUFX3 U567 ( .A(n4321), .Y(n4265) );
  CLKBUFX3 U568 ( .A(n4320), .Y(n4266) );
  CLKBUFX3 U569 ( .A(n4320), .Y(n4267) );
  CLKBUFX3 U570 ( .A(n4320), .Y(n4268) );
  CLKBUFX3 U571 ( .A(n4320), .Y(n4269) );
  CLKBUFX3 U572 ( .A(n4319), .Y(n4270) );
  CLKBUFX3 U573 ( .A(n4319), .Y(n4271) );
  CLKBUFX3 U574 ( .A(n4319), .Y(n4272) );
  CLKBUFX3 U575 ( .A(n4319), .Y(n4273) );
  CLKBUFX3 U576 ( .A(n4318), .Y(n4274) );
  CLKBUFX3 U577 ( .A(n4318), .Y(n4275) );
  CLKBUFX3 U578 ( .A(n4318), .Y(n4276) );
  CLKBUFX3 U579 ( .A(n4318), .Y(n4277) );
  CLKBUFX3 U580 ( .A(n4317), .Y(n4278) );
  CLKBUFX3 U581 ( .A(n4317), .Y(n4279) );
  CLKBUFX3 U582 ( .A(n4317), .Y(n4280) );
  CLKBUFX3 U583 ( .A(n4317), .Y(n4281) );
  CLKBUFX3 U584 ( .A(n4316), .Y(n4282) );
  CLKBUFX3 U585 ( .A(n4316), .Y(n4283) );
  CLKBUFX3 U586 ( .A(n4316), .Y(n4284) );
  CLKBUFX3 U587 ( .A(n4316), .Y(n4285) );
  CLKBUFX3 U588 ( .A(n4315), .Y(n4286) );
  CLKBUFX3 U589 ( .A(n4315), .Y(n4287) );
  CLKBUFX3 U590 ( .A(n4315), .Y(n4288) );
  CLKBUFX3 U591 ( .A(n4315), .Y(n4289) );
  CLKBUFX3 U592 ( .A(n4314), .Y(n4290) );
  CLKBUFX3 U593 ( .A(n4314), .Y(n4291) );
  CLKBUFX3 U594 ( .A(n4314), .Y(n4292) );
  CLKBUFX3 U595 ( .A(n4314), .Y(n4293) );
  CLKBUFX3 U596 ( .A(n4313), .Y(n4294) );
  CLKBUFX3 U597 ( .A(n4313), .Y(n4295) );
  CLKBUFX3 U598 ( .A(n4313), .Y(n4296) );
  CLKBUFX3 U599 ( .A(n4313), .Y(n4297) );
  CLKBUFX3 U600 ( .A(n4312), .Y(n4298) );
  CLKBUFX3 U601 ( .A(n4312), .Y(n4299) );
  CLKBUFX3 U602 ( .A(n4312), .Y(n4300) );
  CLKBUFX3 U603 ( .A(n4312), .Y(n4301) );
  CLKBUFX3 U604 ( .A(n4311), .Y(n4302) );
  CLKBUFX3 U605 ( .A(n4311), .Y(n4303) );
  CLKBUFX3 U606 ( .A(n4311), .Y(n4304) );
  CLKBUFX3 U607 ( .A(n4311), .Y(n4305) );
  CLKBUFX3 U608 ( .A(n4310), .Y(n4306) );
  CLKBUFX3 U609 ( .A(n4310), .Y(n4307) );
  CLKBUFX3 U610 ( .A(n4310), .Y(n4308) );
  CLKBUFX3 U611 ( .A(n4310), .Y(n4309) );
  CLKBUFX3 U612 ( .A(n4335), .Y(n4206) );
  CLKBUFX3 U613 ( .A(n4335), .Y(n4207) );
  CLKBUFX3 U614 ( .A(n4335), .Y(n4208) );
  CLKBUFX3 U615 ( .A(n4335), .Y(n4209) );
  CLKBUFX3 U616 ( .A(n4334), .Y(n4210) );
  CLKBUFX3 U617 ( .A(n4334), .Y(n4211) );
  CLKBUFX3 U618 ( .A(n4334), .Y(n4212) );
  CLKBUFX3 U619 ( .A(n4334), .Y(n4213) );
  CLKBUFX3 U620 ( .A(n4336), .Y(n4333) );
  CLKBUFX3 U621 ( .A(n4336), .Y(n4332) );
  CLKBUFX3 U622 ( .A(n4345), .Y(n4331) );
  CLKBUFX3 U623 ( .A(n4345), .Y(n4330) );
  CLKBUFX3 U624 ( .A(n4337), .Y(n4329) );
  CLKBUFX3 U625 ( .A(n4337), .Y(n4328) );
  CLKBUFX3 U626 ( .A(n4344), .Y(n4327) );
  CLKBUFX3 U627 ( .A(n4344), .Y(n4326) );
  CLKBUFX3 U628 ( .A(n4338), .Y(n4325) );
  CLKBUFX3 U629 ( .A(n4338), .Y(n4324) );
  CLKBUFX3 U630 ( .A(n4343), .Y(n4323) );
  CLKBUFX3 U631 ( .A(n4343), .Y(n4322) );
  CLKBUFX3 U632 ( .A(n4339), .Y(n4321) );
  CLKBUFX3 U633 ( .A(n4339), .Y(n4320) );
  CLKBUFX3 U634 ( .A(n4342), .Y(n4319) );
  CLKBUFX3 U635 ( .A(n4342), .Y(n4318) );
  CLKBUFX3 U636 ( .A(n4341), .Y(n4317) );
  CLKBUFX3 U637 ( .A(n4336), .Y(n4316) );
  CLKBUFX3 U638 ( .A(n4341), .Y(n4315) );
  CLKBUFX3 U639 ( .A(n4337), .Y(n4314) );
  CLKBUFX3 U640 ( .A(n4340), .Y(n4313) );
  CLKBUFX3 U641 ( .A(n4338), .Y(n4312) );
  CLKBUFX3 U642 ( .A(n4340), .Y(n4311) );
  CLKBUFX3 U643 ( .A(n4340), .Y(n4310) );
  CLKBUFX3 U644 ( .A(n1363), .Y(n1546) );
  CLKBUFX3 U645 ( .A(n1359), .Y(n1550) );
  CLKBUFX3 U646 ( .A(n4042), .Y(n4036) );
  CLKBUFX3 U647 ( .A(n4056), .Y(n4050) );
  CLKBUFX3 U648 ( .A(n4090), .Y(n4091) );
  CLKBUFX3 U649 ( .A(n4104), .Y(n4105) );
  CLKBUFX3 U650 ( .A(n4078), .Y(n4080) );
  CLKBUFX3 U651 ( .A(n4184), .Y(n4185) );
  CLKBUFX3 U652 ( .A(n4042), .Y(n4037) );
  CLKBUFX3 U653 ( .A(n4090), .Y(n4092) );
  CLKBUFX3 U654 ( .A(n4104), .Y(n4106) );
  CLKBUFX3 U655 ( .A(n4057), .Y(n4058) );
  CLKBUFX3 U656 ( .A(n4078), .Y(n4081) );
  CLKBUFX3 U657 ( .A(n4184), .Y(n4186) );
  CLKBUFX3 U658 ( .A(n4042), .Y(n4038) );
  CLKBUFX3 U659 ( .A(n4090), .Y(n4093) );
  CLKBUFX3 U660 ( .A(n4104), .Y(n4107) );
  CLKBUFX3 U661 ( .A(n4057), .Y(n4059) );
  CLKBUFX3 U662 ( .A(n4184), .Y(n4187) );
  CLKBUFX3 U663 ( .A(n4042), .Y(n4039) );
  CLKBUFX3 U664 ( .A(n4056), .Y(n4051) );
  CLKBUFX3 U665 ( .A(n4057), .Y(n4060) );
  CLKBUFX3 U666 ( .A(n4184), .Y(n4188) );
  CLKBUFX3 U667 ( .A(n4042), .Y(n4040) );
  CLKBUFX3 U668 ( .A(n1700), .Y(n4052) );
  CLKBUFX3 U669 ( .A(n4104), .Y(n4108) );
  CLKBUFX3 U670 ( .A(n4056), .Y(n4053) );
  CLKBUFX3 U671 ( .A(n4057), .Y(n4061) );
  CLKBUFX3 U672 ( .A(n4056), .Y(n4054) );
  CLKBUFX3 U673 ( .A(n4090), .Y(n4094) );
  CLKBUFX3 U674 ( .A(n4104), .Y(n4109) );
  CLKBUFX3 U675 ( .A(n4057), .Y(n4062) );
  CLKBUFX3 U676 ( .A(n4184), .Y(n4189) );
  CLKBUFX3 U677 ( .A(n4078), .Y(n4082) );
  CLKBUFX3 U678 ( .A(n4042), .Y(n4041) );
  CLKBUFX3 U679 ( .A(n4056), .Y(n4055) );
  CLKBUFX3 U680 ( .A(n4090), .Y(n4095) );
  CLKBUFX3 U681 ( .A(n4104), .Y(n4110) );
  CLKBUFX3 U682 ( .A(n4184), .Y(n4190) );
  CLKBUFX3 U683 ( .A(n4017), .Y(n4018) );
  CLKBUFX3 U684 ( .A(n4017), .Y(n4019) );
  CLKBUFX3 U685 ( .A(n4017), .Y(n4020) );
  CLKBUFX3 U686 ( .A(n4017), .Y(n4021) );
  CLKBUFX3 U687 ( .A(n4090), .Y(n4096) );
  CLKBUFX3 U688 ( .A(n1359), .Y(n1528) );
  CLKBUFX3 U689 ( .A(n1363), .Y(n1370) );
  CLKBUFX3 U690 ( .A(n1359), .Y(n1365) );
  INVX3 U691 ( .A(n1557), .Y(n4149) );
  INVX3 U692 ( .A(n1557), .Y(n4150) );
  INVX3 U693 ( .A(n1556), .Y(n4153) );
  INVX3 U694 ( .A(n1555), .Y(n4156) );
  INVX3 U695 ( .A(n1554), .Y(n4159) );
  INVX3 U696 ( .A(n4165), .Y(n4162) );
  INVX3 U697 ( .A(n4164), .Y(n4163) );
  CLKBUFX3 U698 ( .A(n4345), .Y(n4336) );
  CLKBUFX3 U699 ( .A(n4344), .Y(n4337) );
  CLKBUFX3 U700 ( .A(n4343), .Y(n4338) );
  CLKBUFX3 U701 ( .A(n4342), .Y(n4339) );
  CLKBUFX3 U702 ( .A(n4347), .Y(n4335) );
  CLKBUFX3 U703 ( .A(n4341), .Y(n4334) );
  CLKBUFX3 U704 ( .A(n1358), .Y(n1363) );
  CLKBUFX3 U705 ( .A(n2628), .Y(n3998) );
  CLKBUFX3 U706 ( .A(n1580), .Y(n1701) );
  CLKBUFX3 U707 ( .A(n1704), .Y(n3999) );
  CLKBUFX3 U708 ( .A(n1351), .Y(n1357) );
  INVX3 U709 ( .A(n4120), .Y(n4112) );
  INVX3 U710 ( .A(n4120), .Y(n4118) );
  CLKBUFX3 U711 ( .A(n4078), .Y(n4079) );
  CLKBUFX3 U712 ( .A(n4015), .Y(n4008) );
  CLKBUFX3 U713 ( .A(n4015), .Y(n4009) );
  CLKBUFX3 U714 ( .A(n4015), .Y(n4010) );
  CLKBUFX3 U715 ( .A(n4015), .Y(n4011) );
  CLKBUFX3 U716 ( .A(n4015), .Y(n4012) );
  CLKBUFX3 U717 ( .A(n4015), .Y(n4013) );
  CLKBUFX3 U718 ( .A(n4015), .Y(n4014) );
  CLKBUFX3 U719 ( .A(n1693), .Y(n1697) );
  CLKBUFX3 U720 ( .A(n1704), .Y(n3997) );
  CLKBUFX3 U721 ( .A(n3997), .Y(n3996) );
  CLKBUFX3 U722 ( .A(n1693), .Y(n1696) );
  CLKBUFX3 U723 ( .A(n3998), .Y(n3995) );
  CLKBUFX3 U724 ( .A(n1693), .Y(n1695) );
  CLKBUFX3 U725 ( .A(n1351), .Y(n1355) );
  CLKBUFX3 U726 ( .A(n1351), .Y(n1356) );
  INVX3 U727 ( .A(n4119), .Y(n4117) );
  INVX3 U728 ( .A(n4120), .Y(n4116) );
  INVX3 U729 ( .A(n4120), .Y(n4113) );
  INVX3 U730 ( .A(n4119), .Y(n4115) );
  INVX3 U731 ( .A(n4119), .Y(n4114) );
  CLKBUFX3 U732 ( .A(n4071), .Y(n4076) );
  CLKBUFX3 U733 ( .A(n8), .Y(n4068) );
  CLKBUFX3 U734 ( .A(n4071), .Y(n4075) );
  CLKBUFX3 U735 ( .A(n8), .Y(n4067) );
  CLKBUFX3 U736 ( .A(n8), .Y(n4065) );
  CLKBUFX3 U737 ( .A(n8), .Y(n4066) );
  CLKBUFX3 U738 ( .A(n4071), .Y(n4073) );
  CLKBUFX3 U739 ( .A(n4071), .Y(n4074) );
  CLKBUFX3 U740 ( .A(n4065), .Y(n4070) );
  CLKBUFX3 U741 ( .A(n4066), .Y(n4069) );
  CLKBUFX3 U742 ( .A(n1554), .Y(n4160) );
  CLKBUFX3 U743 ( .A(n11), .Y(n4164) );
  CLKBUFX3 U744 ( .A(n11), .Y(n4165) );
  CLKBUFX3 U745 ( .A(n6), .Y(n4023) );
  CLKBUFX3 U746 ( .A(n6), .Y(n4024) );
  CLKBUFX3 U747 ( .A(n4027), .Y(n4025) );
  CLKBUFX3 U748 ( .A(n4027), .Y(n4026) );
  CLKBUFX3 U749 ( .A(n6), .Y(n4027) );
  CLKBUFX3 U750 ( .A(n6), .Y(n4028) );
  CLKBUFX3 U751 ( .A(n6), .Y(n4022) );
  CLKBUFX3 U752 ( .A(n4049), .Y(n4044) );
  CLKBUFX3 U753 ( .A(n4088), .Y(n4085) );
  CLKBUFX3 U754 ( .A(n4097), .Y(n4099) );
  CLKBUFX3 U755 ( .A(n2), .Y(n4178) );
  CLKBUFX3 U756 ( .A(n4035), .Y(n4030) );
  CLKBUFX3 U757 ( .A(n4049), .Y(n4045) );
  CLKBUFX3 U758 ( .A(n4098), .Y(n4100) );
  CLKBUFX3 U759 ( .A(n2), .Y(n4179) );
  CLKBUFX3 U760 ( .A(n4035), .Y(n4031) );
  CLKBUFX3 U761 ( .A(n4049), .Y(n4046) );
  CLKBUFX3 U762 ( .A(n7), .Y(n4086) );
  CLKBUFX3 U763 ( .A(n4181), .Y(n4180) );
  CLKBUFX3 U764 ( .A(n4035), .Y(n4032) );
  CLKBUFX3 U765 ( .A(n4049), .Y(n4047) );
  CLKBUFX3 U766 ( .A(n4098), .Y(n4101) );
  CLKBUFX3 U767 ( .A(n4035), .Y(n4033) );
  CLKBUFX3 U768 ( .A(n7), .Y(n4087) );
  CLKBUFX3 U769 ( .A(n7), .Y(n4088) );
  CLKBUFX3 U770 ( .A(n5), .Y(n4102) );
  CLKBUFX3 U771 ( .A(n2), .Y(n4181) );
  CLKBUFX3 U772 ( .A(n4035), .Y(n4034) );
  CLKBUFX3 U773 ( .A(n4049), .Y(n4048) );
  CLKBUFX3 U774 ( .A(n7), .Y(n4089) );
  CLKBUFX3 U775 ( .A(n5), .Y(n4103) );
  CLKBUFX3 U776 ( .A(n4181), .Y(n4182) );
  CLKBUFX3 U777 ( .A(n2), .Y(n4183) );
  CLKBUFX3 U778 ( .A(n4035), .Y(n4029) );
  CLKBUFX3 U779 ( .A(n4049), .Y(n4043) );
  CLKBUFX3 U780 ( .A(n4071), .Y(n4077) );
  CLKBUFX3 U781 ( .A(n7), .Y(n4084) );
  CLKBUFX3 U782 ( .A(n5), .Y(n4098) );
  INVX3 U783 ( .A(n4175), .Y(n4174) );
  INVX3 U784 ( .A(n4169), .Y(n4166) );
  INVX3 U785 ( .A(n4168), .Y(n4167) );
  INVX3 U786 ( .A(n1547), .Y(n4170) );
  INVX3 U787 ( .A(n4176), .Y(n4173) );
  CLKBUFX3 U788 ( .A(n1557), .Y(n4151) );
  CLKBUFX3 U789 ( .A(n1556), .Y(n4154) );
  CLKBUFX3 U790 ( .A(n1555), .Y(n4157) );
  CLKBUFX3 U791 ( .A(n1554), .Y(n4161) );
  CLKBUFX3 U792 ( .A(n1344), .Y(n1348) );
  CLKBUFX3 U793 ( .A(n1343), .Y(n1347) );
  CLKBUFX3 U794 ( .A(n1344), .Y(n1346) );
  CLKBUFX3 U795 ( .A(n1343), .Y(n1345) );
  CLKBUFX3 U796 ( .A(n1349), .Y(n1344) );
  CLKBUFX3 U797 ( .A(mem_read), .Y(n1343) );
  CLKBUFX3 U798 ( .A(n4347), .Y(n4341) );
  CLKBUFX3 U799 ( .A(n4347), .Y(n4340) );
  CLKBUFX3 U800 ( .A(n4346), .Y(n4345) );
  CLKBUFX3 U801 ( .A(n4346), .Y(n4344) );
  CLKBUFX3 U802 ( .A(n4346), .Y(n4343) );
  CLKBUFX3 U803 ( .A(n4346), .Y(n4342) );
  CLKBUFX3 U804 ( .A(n1552), .Y(n1580) );
  CLKBUFX3 U805 ( .A(n1350), .Y(n1353) );
  INVX3 U806 ( .A(n4140), .Y(n4132) );
  INVX3 U807 ( .A(n4130), .Y(n4122) );
  CLKBUFX3 U808 ( .A(n1359), .Y(n1358) );
  CLKBUFX3 U809 ( .A(n4357), .Y(n1359) );
  CLKBUFX3 U810 ( .A(n1703), .Y(n2628) );
  INVX3 U811 ( .A(n1299), .Y(n4141) );
  INVX3 U812 ( .A(n4139), .Y(n4137) );
  INVX3 U813 ( .A(n4139), .Y(n4138) );
  INVX3 U814 ( .A(n4129), .Y(n4127) );
  INVX3 U815 ( .A(n1299), .Y(n4147) );
  INVX3 U816 ( .A(n4129), .Y(n4128) );
  INVX3 U817 ( .A(n1299), .Y(n4148) );
  CLKBUFX3 U818 ( .A(n4015), .Y(n4007) );
  CLKBUFX3 U819 ( .A(n1707), .Y(n4015) );
  CLKBUFX3 U820 ( .A(n1694), .Y(n4078) );
  CLKBUFX3 U821 ( .A(n1692), .Y(n4090) );
  CLKBUFX3 U822 ( .A(n1578), .Y(n4104) );
  CLKBUFX3 U823 ( .A(n1705), .Y(n4017) );
  CLKBUFX3 U824 ( .A(n1702), .Y(n4042) );
  CLKBUFX3 U825 ( .A(n1700), .Y(n4056) );
  CLKBUFX3 U826 ( .A(n1552), .Y(n1693) );
  CLKBUFX3 U827 ( .A(n1350), .Y(n1354) );
  INVX3 U828 ( .A(n4139), .Y(n4136) );
  INVX3 U829 ( .A(n4140), .Y(n4133) );
  INVX3 U830 ( .A(n4139), .Y(n4135) );
  INVX3 U831 ( .A(n4139), .Y(n4134) );
  INVX3 U832 ( .A(n1299), .Y(n4145) );
  INVX3 U833 ( .A(n4129), .Y(n4126) );
  INVX3 U834 ( .A(n1299), .Y(n4146) );
  INVX3 U835 ( .A(n1299), .Y(n4144) );
  INVX3 U836 ( .A(n4130), .Y(n4123) );
  INVX3 U837 ( .A(n4129), .Y(n4125) );
  INVX3 U838 ( .A(n1299), .Y(n4143) );
  INVX3 U839 ( .A(n4129), .Y(n4124) );
  INVX3 U840 ( .A(n1299), .Y(n4142) );
  CLKBUFX3 U841 ( .A(n1368), .Y(n4196) );
  CLKBUFX3 U842 ( .A(n1728), .Y(n4005) );
  CLKBUFX3 U843 ( .A(n1795), .Y(n4003) );
  CLKBUFX3 U844 ( .A(n1761), .Y(n4004) );
  CLKBUFX3 U845 ( .A(n1709), .Y(n4006) );
  INVX4 U846 ( .A(n4001), .Y(n4000) );
  CLKBUFX3 U847 ( .A(n4071), .Y(n4072) );
  CLKBUFX3 U848 ( .A(n13), .Y(n4175) );
  CLKBUFX3 U849 ( .A(n13), .Y(n4176) );
  CLKBUFX3 U850 ( .A(n12), .Y(n4168) );
  CLKBUFX3 U851 ( .A(n12), .Y(n4169) );
  CLKBUFX3 U852 ( .A(n4194), .Y(n4195) );
  CLKBUFX3 U853 ( .A(n8), .Y(n4064) );
  CLKBUFX3 U854 ( .A(n2), .Y(n4177) );
  CLKBUFX3 U855 ( .A(n7), .Y(n4083) );
  CLKBUFX3 U856 ( .A(n5), .Y(n4097) );
  CLKBUFX3 U857 ( .A(n1547), .Y(n4171) );
  CLKBUFX3 U858 ( .A(n1341), .Y(n1349) );
  CLKBUFX3 U859 ( .A(n1342), .Y(n1341) );
  CLKBUFX3 U860 ( .A(n1556), .Y(n4155) );
  CLKBUFX3 U861 ( .A(n1555), .Y(n4158) );
  CLKBUFX3 U862 ( .A(n1557), .Y(n4152) );
  CLKBUFX3 U863 ( .A(n3), .Y(n4035) );
  CLKBUFX3 U864 ( .A(n4), .Y(n4049) );
  CLKBUFX3 U865 ( .A(n4120), .Y(n4119) );
  CLKINVX1 U866 ( .A(n4205), .Y(n4347) );
  CLKINVX1 U867 ( .A(n1553), .Y(n4357) );
  CLKBUFX3 U868 ( .A(n1352), .Y(n1350) );
  CLKBUFX3 U869 ( .A(n4356), .Y(n1352) );
  CLKBUFX3 U870 ( .A(n1558), .Y(n1552) );
  CLKBUFX3 U871 ( .A(n4359), .Y(n1558) );
  NOR2BX1 U872 ( .AN(n1691), .B(n4116), .Y(n1699) );
  NOR2BX1 U873 ( .AN(n1691), .B(n4128), .Y(n1694) );
  NOR2BX1 U874 ( .AN(n1691), .B(n4133), .Y(n1692) );
  NOR2BX1 U875 ( .AN(n1691), .B(n4145), .Y(n1578) );
  NOR2BX1 U876 ( .AN(n1691), .B(n1354), .Y(n1705) );
  NOR2BX1 U877 ( .AN(n1691), .B(n1552), .Y(n1702) );
  NOR2BX1 U878 ( .AN(n1691), .B(n1528), .Y(n1700) );
  CLKBUFX3 U879 ( .A(n1526), .Y(n4184) );
  NOR2BX1 U880 ( .AN(n1691), .B(n3999), .Y(n1526) );
  CLKBUFX3 U881 ( .A(n4140), .Y(n4139) );
  CLKBUFX3 U882 ( .A(n4356), .Y(n1351) );
  CLKBUFX3 U883 ( .A(n1704), .Y(n1703) );
  CLKBUFX3 U884 ( .A(n4360), .Y(n1704) );
  CLKINVX1 U885 ( .A(n4111), .Y(n4120) );
  AND3X2 U886 ( .A(n4200), .B(n4194), .C(n4204), .Y(n1728) );
  AND3X2 U887 ( .A(n4200), .B(n4193), .C(n4204), .Y(n1709) );
  AND2X2 U888 ( .A(n1793), .B(n4204), .Y(n1795) );
  AND2X2 U889 ( .A(n1793), .B(n4200), .Y(n1761) );
  CLKBUFX3 U890 ( .A(n1706), .Y(n4016) );
  CLKBUFX3 U891 ( .A(n1698), .Y(n4063) );
  CLKBUFX3 U892 ( .A(n14), .Y(n4001) );
  CLKBUFX3 U893 ( .A(n14), .Y(n4002) );
  INVX3 U894 ( .A(n1294), .Y(n1338) );
  INVX3 U895 ( .A(n1294), .Y(n1339) );
  AND2X2 U896 ( .A(n4193), .B(n4196), .Y(n1793) );
  CLKBUFX3 U897 ( .A(n1368), .Y(n4194) );
  NAND2X1 U898 ( .A(n1548), .B(n1299), .Y(n1557) );
  CLKINVX1 U899 ( .A(n1565), .Y(n4349) );
  CLKBUFX3 U900 ( .A(n4197), .Y(n4198) );
  CLKBUFX3 U901 ( .A(n4204), .Y(n4203) );
  CLKBUFX3 U902 ( .A(n4200), .Y(n4199) );
  CLKBUFX3 U903 ( .A(n4201), .Y(n4202) );
  CLKBUFX3 U904 ( .A(n4193), .Y(n4192) );
  CLKBUFX3 U905 ( .A(n1547), .Y(n4172) );
  CLKBUFX3 U906 ( .A(n4348), .Y(n1342) );
  CLKBUFX3 U907 ( .A(n1), .Y(n4071) );
  AND2X2 U908 ( .A(n1548), .B(n4139), .Y(n1295) );
  CLKINVX1 U909 ( .A(n1295), .Y(n1556) );
  AND2X2 U910 ( .A(n1548), .B(n4129), .Y(n1296) );
  CLKINVX1 U911 ( .A(n1296), .Y(n1555) );
  AND2X2 U912 ( .A(n1548), .B(n4119), .Y(n1297) );
  CLKINVX1 U913 ( .A(n1297), .Y(n1554) );
  CLKBUFX3 U914 ( .A(n4130), .Y(n4129) );
  CLKBUFX3 U915 ( .A(proc_reset), .Y(n4205) );
  NOR3X1 U916 ( .A(n4358), .B(mem_addr[2]), .C(n4361), .Y(n1553) );
  NOR4X1 U917 ( .A(n2016), .B(n2017), .C(n2018), .D(n2019), .Y(n1981) );
  NAND4X1 U918 ( .A(n2020), .B(n2021), .C(n2022), .D(n2023), .Y(n2019) );
  NAND4X1 U919 ( .A(n2035), .B(n2036), .C(n2037), .D(n2038), .Y(n2017) );
  NAND4X1 U920 ( .A(n2027), .B(n2028), .C(n2029), .D(n2030), .Y(n2018) );
  NOR4X1 U921 ( .A(n1880), .B(n1881), .C(n1882), .D(n1883), .Y(n1845) );
  NAND4X1 U922 ( .A(n1884), .B(n1885), .C(n1886), .D(n1887), .Y(n1883) );
  NAND4X1 U923 ( .A(n1899), .B(n1900), .C(n1901), .D(n1902), .Y(n1881) );
  NAND4X1 U924 ( .A(n1891), .B(n1892), .C(n1893), .D(n1894), .Y(n1882) );
  NOR4X1 U925 ( .A(n2082), .B(n2083), .C(n2084), .D(n2085), .Y(n1979) );
  NAND4X1 U926 ( .A(n2086), .B(n2087), .C(n2088), .D(n2089), .Y(n2085) );
  NAND4X1 U927 ( .A(n2101), .B(n2102), .C(n2103), .D(n2104), .Y(n2083) );
  NAND4X1 U928 ( .A(n2093), .B(n2094), .C(n2095), .D(n2096), .Y(n2084) );
  NOR4X1 U929 ( .A(n2049), .B(n2050), .C(n2051), .D(n2052), .Y(n1980) );
  NAND4X1 U930 ( .A(n2053), .B(n2054), .C(n2055), .D(n2056), .Y(n2052) );
  NAND4X1 U931 ( .A(n2068), .B(n2069), .C(n2070), .D(n2071), .Y(n2050) );
  NAND4X1 U932 ( .A(n2060), .B(n2061), .C(n2062), .D(n2063), .Y(n2051) );
  NOR4X1 U933 ( .A(n1913), .B(n1914), .C(n1915), .D(n1916), .Y(n1844) );
  NAND4X1 U934 ( .A(n1917), .B(n1918), .C(n1919), .D(n1920), .Y(n1916) );
  NAND4X1 U935 ( .A(n1932), .B(n1933), .C(n1934), .D(n1935), .Y(n1914) );
  NAND4X1 U936 ( .A(n1924), .B(n1925), .C(n1926), .D(n1927), .Y(n1915) );
  CLKINVX1 U937 ( .A(n1549), .Y(n4356) );
  CLKINVX1 U938 ( .A(n1551), .Y(n4359) );
  AND2X2 U939 ( .A(n1841), .B(n1842), .Y(n1569) );
  NOR4X1 U940 ( .A(n1843), .B(n1844), .C(n1845), .D(n1846), .Y(n1842) );
  NOR4X1 U941 ( .A(n1979), .B(n1980), .C(n1981), .D(n1982), .Y(n1841) );
  NOR4X1 U942 ( .A(n1847), .B(n1848), .C(n1849), .D(n1850), .Y(n1846) );
  CLKINVX1 U943 ( .A(n4121), .Y(n4130) );
  CLKINVX1 U944 ( .A(n4131), .Y(n4140) );
  NOR2BX1 U945 ( .AN(n1575), .B(n1569), .Y(n1707) );
  NAND2X1 U946 ( .A(n1575), .B(n1569), .Y(n1570) );
  NOR4X1 U947 ( .A(n1983), .B(n1984), .C(n1985), .D(n1986), .Y(n1982) );
  NAND4X1 U948 ( .A(n2010), .B(n2011), .C(n2012), .D(n2013), .Y(n1983) );
  NAND4X1 U949 ( .A(n1987), .B(n1988), .C(n1989), .D(n1990), .Y(n1986) );
  NAND4X1 U950 ( .A(n2002), .B(n2003), .C(n2004), .D(n2005), .Y(n1984) );
  NOR4X1 U951 ( .A(n1946), .B(n1947), .C(n1948), .D(n1949), .Y(n1843) );
  NAND4X1 U952 ( .A(n1950), .B(n1951), .C(n1952), .D(n1953), .Y(n1949) );
  NAND4X1 U953 ( .A(n1965), .B(n1966), .C(n1967), .D(n1968), .Y(n1947) );
  NAND4X1 U954 ( .A(n1957), .B(n1958), .C(n1959), .D(n1960), .Y(n1948) );
  CLKINVX1 U955 ( .A(n1577), .Y(n4360) );
  AND2X2 U956 ( .A(n1570), .B(n1337), .Y(n1691) );
  CLKBUFX3 U957 ( .A(n1562), .Y(n4111) );
  NAND3X1 U958 ( .A(n4358), .B(n4361), .C(mem_addr[2]), .Y(n1562) );
  NAND2X1 U959 ( .A(n4354), .B(n4355), .Y(n1368) );
  AND3X2 U960 ( .A(n1570), .B(n1549), .C(n1337), .Y(n1706) );
  AND3X2 U961 ( .A(n1570), .B(n4119), .C(n1337), .Y(n1698) );
  CLKBUFX3 U962 ( .A(n4197), .Y(n4200) );
  CLKBUFX3 U963 ( .A(n10), .Y(n4197) );
  CLKBUFX3 U964 ( .A(n4201), .Y(n4204) );
  CLKBUFX3 U965 ( .A(n9), .Y(n4201) );
  OAI21X1 U966 ( .A0(n1575), .A1(n4418), .B0(n1340), .Y(n1565) );
  CLKINVX1 U967 ( .A(n1361), .Y(n4348) );
  CLKBUFX3 U968 ( .A(n4191), .Y(n4193) );
  CLKBUFX3 U969 ( .A(n16), .Y(n4191) );
  AND2X2 U970 ( .A(n1548), .B(n1549), .Y(n1298) );
  CLKINVX1 U971 ( .A(n1298), .Y(n1547) );
  INVX1 U972 ( .A(proc_addr[3]), .Y(n4361) );
  INVX1 U973 ( .A(proc_addr[2]), .Y(n4358) );
  CLKBUFX3 U974 ( .A(n1561), .Y(n4121) );
  NAND3XL U975 ( .A(proc_addr[2]), .B(n4361), .C(mem_addr[2]), .Y(n1561) );
  INVX16 U976 ( .A(n1335), .Y(mem_addr[2]) );
  NOR4X1 U977 ( .A(n1353), .B(n49), .C(n2047), .D(n2048), .Y(n2046) );
  XOR2XL U978 ( .A(\tag_r[1][4] ), .B(proc_addr[9]), .Y(n2047) );
  XOR2XL U979 ( .A(\tag_r[1][6] ), .B(proc_addr[11]), .Y(n2048) );
  NOR4X1 U980 ( .A(n1580), .B(n48), .C(n2080), .D(n2081), .Y(n2079) );
  XOR2XL U981 ( .A(\tag_r[2][4] ), .B(proc_addr[9]), .Y(n2080) );
  XOR2XL U982 ( .A(\tag_r[2][6] ), .B(proc_addr[11]), .Y(n2081) );
  NOR4X1 U983 ( .A(n1363), .B(n47), .C(n2113), .D(n2114), .Y(n2112) );
  XOR2XL U984 ( .A(\tag_r[3][4] ), .B(proc_addr[9]), .Y(n2113) );
  XOR2XL U985 ( .A(\tag_r[3][6] ), .B(proc_addr[11]), .Y(n2114) );
  NOR4X1 U986 ( .A(n4122), .B(n45), .C(n1911), .D(n1912), .Y(n1910) );
  XOR2XL U987 ( .A(\tag_r[5][4] ), .B(proc_addr[9]), .Y(n1911) );
  XOR2XL U988 ( .A(\tag_r[5][6] ), .B(proc_addr[11]), .Y(n1912) );
  NOR4X1 U989 ( .A(n4132), .B(n44), .C(n1944), .D(n1945), .Y(n1943) );
  XOR2XL U990 ( .A(\tag_r[6][4] ), .B(proc_addr[9]), .Y(n1944) );
  XOR2XL U991 ( .A(\tag_r[6][6] ), .B(proc_addr[11]), .Y(n1945) );
  NAND4X1 U992 ( .A(n2043), .B(n2044), .C(n2045), .D(n2046), .Y(n2016) );
  XOR2XL U993 ( .A(n1253), .B(proc_addr[15]), .Y(n2045) );
  XOR2XL U994 ( .A(n1258), .B(proc_addr[10]), .Y(n2044) );
  XOR2XL U995 ( .A(n1252), .B(proc_addr[16]), .Y(n2043) );
  NAND4X1 U996 ( .A(n2076), .B(n2077), .C(n2078), .D(n2079), .Y(n2049) );
  XOR2XL U997 ( .A(n1228), .B(proc_addr[15]), .Y(n2078) );
  XOR2XL U998 ( .A(n1233), .B(proc_addr[10]), .Y(n2077) );
  XOR2XL U999 ( .A(n1227), .B(proc_addr[16]), .Y(n2076) );
  NAND4X1 U1000 ( .A(n2109), .B(n2110), .C(n2111), .D(n2112), .Y(n2082) );
  XOR2XL U1001 ( .A(n1203), .B(proc_addr[15]), .Y(n2111) );
  XOR2XL U1002 ( .A(n1208), .B(proc_addr[10]), .Y(n2110) );
  XOR2XL U1003 ( .A(n1202), .B(proc_addr[16]), .Y(n2109) );
  NAND4X1 U1004 ( .A(n1907), .B(n1908), .C(n1909), .D(n1910), .Y(n1880) );
  XOR2XL U1005 ( .A(n1153), .B(proc_addr[15]), .Y(n1909) );
  XOR2XL U1006 ( .A(n1158), .B(proc_addr[10]), .Y(n1908) );
  XOR2XL U1007 ( .A(n1152), .B(proc_addr[16]), .Y(n1907) );
  NAND4X1 U1008 ( .A(n1940), .B(n1941), .C(n1942), .D(n1943), .Y(n1913) );
  XOR2XL U1009 ( .A(n1128), .B(proc_addr[15]), .Y(n1942) );
  XOR2XL U1010 ( .A(n1133), .B(proc_addr[10]), .Y(n1941) );
  XOR2XL U1011 ( .A(n1127), .B(proc_addr[16]), .Y(n1940) );
  NAND3X1 U1012 ( .A(n1568), .B(n64), .C(n1569), .Y(n1360) );
  NAND3X1 U1013 ( .A(n1360), .B(n61), .C(n1361), .Y(proc_stall) );
  CLKBUFX3 U1014 ( .A(n1560), .Y(n4131) );
  NAND3XL U1015 ( .A(proc_addr[3]), .B(n4358), .C(mem_addr[2]), .Y(n1560) );
  NOR4X1 U1016 ( .A(n2659), .B(n2660), .C(n2661), .D(n2662), .Y(n2658) );
  OAI22XL U1017 ( .A0(n4138), .A1(n1138), .B0(n4148), .B1(n1113), .Y(n2659) );
  OAI22XL U1018 ( .A0(n4113), .A1(n1188), .B0(n4128), .B1(n1163), .Y(n2660) );
  NOR4X1 U1019 ( .A(n2654), .B(n2655), .C(n2656), .D(n2657), .Y(n2653) );
  OAI22XL U1020 ( .A0(n4138), .A1(n1137), .B0(n4148), .B1(n1112), .Y(n2654) );
  OAI22XL U1021 ( .A0(n4113), .A1(n1187), .B0(n4128), .B1(n1162), .Y(n2655) );
  NOR4X1 U1022 ( .A(n2649), .B(n2650), .C(n2651), .D(n2652), .Y(n2648) );
  OAI22XL U1023 ( .A0(n4138), .A1(n1136), .B0(n4148), .B1(n1111), .Y(n2649) );
  OAI22XL U1024 ( .A0(n4118), .A1(n1186), .B0(n4128), .B1(n1161), .Y(n2650) );
  NOR4X1 U1025 ( .A(n2644), .B(n2645), .C(n2646), .D(n2647), .Y(n2643) );
  OAI22XL U1026 ( .A0(n4138), .A1(n1135), .B0(n4148), .B1(n1110), .Y(n2644) );
  OAI22XL U1027 ( .A0(n4118), .A1(n1185), .B0(n4128), .B1(n1160), .Y(n2645) );
  NOR4X1 U1028 ( .A(n2639), .B(n2640), .C(n2641), .D(n2642), .Y(n2638) );
  OAI22XL U1029 ( .A0(n4137), .A1(n1134), .B0(n4147), .B1(n1109), .Y(n2639) );
  OAI22XL U1030 ( .A0(n4118), .A1(n1184), .B0(n4127), .B1(n1159), .Y(n2640) );
  NOR4X1 U1031 ( .A(n2634), .B(n2635), .C(n2636), .D(n2637), .Y(n2633) );
  OAI22XL U1032 ( .A0(n4137), .A1(n1133), .B0(n4147), .B1(n1108), .Y(n2634) );
  OAI22XL U1033 ( .A0(n4118), .A1(n1183), .B0(n4127), .B1(n1158), .Y(n2635) );
  NOR4X1 U1034 ( .A(n2629), .B(n2630), .C(n2631), .D(n2632), .Y(n2627) );
  OAI22XL U1035 ( .A0(n4137), .A1(n1132), .B0(n4147), .B1(n1107), .Y(n2629) );
  NOR4X1 U1036 ( .A(n2749), .B(n2750), .C(n2751), .D(n2752), .Y(n2748) );
  OAI22XL U1037 ( .A0(n4132), .A1(n1131), .B0(n4141), .B1(n1106), .Y(n2749) );
  OAI22XL U1038 ( .A0(n4112), .A1(n1181), .B0(n4122), .B1(n1156), .Y(n2750) );
  NOR4X1 U1039 ( .A(n2744), .B(n2745), .C(n2746), .D(n2747), .Y(n2743) );
  OAI22XL U1040 ( .A0(n4138), .A1(n1130), .B0(n4145), .B1(n1105), .Y(n2744) );
  OAI22XL U1041 ( .A0(n4118), .A1(n1180), .B0(n4128), .B1(n1155), .Y(n2745) );
  NOR4X1 U1042 ( .A(n2739), .B(n2740), .C(n2741), .D(n2742), .Y(n2738) );
  OAI22XL U1043 ( .A0(n4138), .A1(n1129), .B0(n4143), .B1(n1104), .Y(n2739) );
  OAI22XL U1044 ( .A0(n4117), .A1(n1179), .B0(n4128), .B1(n1154), .Y(n2740) );
  NOR4X1 U1045 ( .A(n2734), .B(n2735), .C(n2736), .D(n2737), .Y(n2733) );
  OAI22XL U1046 ( .A0(n4138), .A1(n1128), .B0(n4142), .B1(n1103), .Y(n2734) );
  OAI22XL U1047 ( .A0(n4118), .A1(n1178), .B0(n4128), .B1(n1153), .Y(n2735) );
  NOR4X1 U1048 ( .A(n2729), .B(n2730), .C(n2731), .D(n2732), .Y(n2728) );
  OAI22XL U1049 ( .A0(n4138), .A1(n1127), .B0(n4144), .B1(n1102), .Y(n2729) );
  OAI22XL U1050 ( .A0(n4117), .A1(n1177), .B0(n4123), .B1(n1152), .Y(n2730) );
  NOR4X1 U1051 ( .A(n2724), .B(n2725), .C(n2726), .D(n2727), .Y(n2723) );
  OAI22XL U1052 ( .A0(n4138), .A1(n1126), .B0(n4148), .B1(n1101), .Y(n2724) );
  OAI22XL U1053 ( .A0(n4117), .A1(n1176), .B0(n4128), .B1(n1151), .Y(n2725) );
  NOR4X1 U1054 ( .A(n2719), .B(n2720), .C(n2721), .D(n2722), .Y(n2718) );
  OAI22XL U1055 ( .A0(n4138), .A1(n1125), .B0(n4148), .B1(n1100), .Y(n2719) );
  OAI22XL U1056 ( .A0(n4113), .A1(n1175), .B0(n4128), .B1(n1150), .Y(n2720) );
  NOR4X1 U1057 ( .A(n2714), .B(n2715), .C(n2716), .D(n2717), .Y(n2713) );
  OAI22XL U1058 ( .A0(n4138), .A1(n1124), .B0(n4148), .B1(n1099), .Y(n2714) );
  OAI22XL U1059 ( .A0(n4115), .A1(n1174), .B0(n4128), .B1(n1149), .Y(n2715) );
  NOR4X1 U1060 ( .A(n2709), .B(n2710), .C(n2711), .D(n2712), .Y(n2708) );
  OAI22XL U1061 ( .A0(n4138), .A1(n1123), .B0(n4148), .B1(n1098), .Y(n2709) );
  OAI22XL U1062 ( .A0(n4114), .A1(n1173), .B0(n4128), .B1(n1148), .Y(n2710) );
  NOR4X1 U1063 ( .A(n2704), .B(n2705), .C(n2706), .D(n2707), .Y(n2703) );
  OAI22XL U1064 ( .A0(n4138), .A1(n1122), .B0(n4148), .B1(n1097), .Y(n2704) );
  OAI22XL U1065 ( .A0(n4111), .A1(n1172), .B0(n4128), .B1(n1147), .Y(n2705) );
  NOR4X1 U1066 ( .A(n2699), .B(n2700), .C(n2701), .D(n2702), .Y(n2698) );
  OAI22XL U1067 ( .A0(n4138), .A1(n1121), .B0(n4148), .B1(n1096), .Y(n2699) );
  OAI22XL U1068 ( .A0(n4115), .A1(n1171), .B0(n4128), .B1(n1146), .Y(n2700) );
  NOR4X1 U1069 ( .A(n2694), .B(n2695), .C(n2696), .D(n2697), .Y(n2693) );
  OAI22XL U1070 ( .A0(n4138), .A1(n1120), .B0(n4148), .B1(n1095), .Y(n2694) );
  OAI22XL U1071 ( .A0(n4117), .A1(n1170), .B0(n4128), .B1(n1145), .Y(n2695) );
  NOR4X1 U1072 ( .A(n2689), .B(n2690), .C(n2691), .D(n2692), .Y(n2688) );
  OAI22XL U1073 ( .A0(n4138), .A1(n1119), .B0(n4148), .B1(n1094), .Y(n2689) );
  OAI22XL U1074 ( .A0(n4114), .A1(n1169), .B0(n4128), .B1(n1144), .Y(n2690) );
  NOR4X1 U1075 ( .A(n2684), .B(n2685), .C(n2686), .D(n2687), .Y(n2683) );
  OAI22XL U1076 ( .A0(n4138), .A1(n1118), .B0(n4148), .B1(n1093), .Y(n2684) );
  OAI22XL U1077 ( .A0(n4116), .A1(n1168), .B0(n4128), .B1(n1143), .Y(n2685) );
  NOR4X1 U1078 ( .A(n2679), .B(n2680), .C(n2681), .D(n2682), .Y(n2678) );
  OAI22XL U1079 ( .A0(n4138), .A1(n1117), .B0(n4148), .B1(n1092), .Y(n2679) );
  OAI22XL U1080 ( .A0(n4113), .A1(n1167), .B0(n4128), .B1(n1142), .Y(n2680) );
  NOR4X1 U1081 ( .A(n2674), .B(n2675), .C(n2676), .D(n2677), .Y(n2673) );
  OAI22XL U1082 ( .A0(n4138), .A1(n1116), .B0(n4148), .B1(n1091), .Y(n2674) );
  OAI22XL U1083 ( .A0(n4111), .A1(n1166), .B0(n4128), .B1(n1141), .Y(n2675) );
  NOR4X1 U1084 ( .A(n2669), .B(n2670), .C(n2671), .D(n2672), .Y(n2668) );
  OAI22XL U1085 ( .A0(n4138), .A1(n1115), .B0(n4148), .B1(n1090), .Y(n2669) );
  OAI22XL U1086 ( .A0(n4115), .A1(n1165), .B0(n4128), .B1(n1140), .Y(n2670) );
  NOR4X1 U1087 ( .A(n2664), .B(n2665), .C(n2666), .D(n2667), .Y(n2663) );
  OAI22XL U1088 ( .A0(n4138), .A1(n1114), .B0(n4148), .B1(n1089), .Y(n2664) );
  OAI22XL U1089 ( .A0(n4114), .A1(n1164), .B0(n4128), .B1(n1139), .Y(n2665) );
  AOI22X2 U1090 ( .A0(mem_rdata[19]), .A1(n1349), .B0(n4007), .B1(n1839), .Y(
        n1688) );
  OAI22XL U1091 ( .A0(n4196), .A1(n4404), .B0(n1474), .B1(n4006), .Y(n1839) );
  AOI22X2 U1092 ( .A0(mem_rdata[20]), .A1(n1349), .B0(n4007), .B1(n1838), .Y(
        n1687) );
  OAI22XL U1093 ( .A0(n4196), .A1(n4405), .B0(n1464), .B1(n4006), .Y(n1838) );
  AOI22X2 U1094 ( .A0(mem_rdata[21]), .A1(n1349), .B0(n4007), .B1(n1837), .Y(
        n1686) );
  OAI22XL U1095 ( .A0(n4196), .A1(n4406), .B0(n1459), .B1(n4006), .Y(n1837) );
  AOI22X2 U1096 ( .A0(mem_rdata[22]), .A1(n1349), .B0(n4007), .B1(n1836), .Y(
        n1685) );
  OAI22XL U1097 ( .A0(n4196), .A1(n4407), .B0(n1454), .B1(n4006), .Y(n1836) );
  AOI22X2 U1098 ( .A0(mem_rdata[23]), .A1(n1349), .B0(n4007), .B1(n1835), .Y(
        n1684) );
  OAI22XL U1099 ( .A0(n4195), .A1(n4408), .B0(n1449), .B1(n4006), .Y(n1835) );
  AOI22X2 U1100 ( .A0(mem_rdata[24]), .A1(n1349), .B0(n4007), .B1(n1834), .Y(
        n1683) );
  OAI22XL U1101 ( .A0(n4196), .A1(n4409), .B0(n1444), .B1(n4006), .Y(n1834) );
  AOI22X2 U1102 ( .A0(mem_rdata[25]), .A1(n1349), .B0(n4007), .B1(n1833), .Y(
        n1682) );
  OAI22XL U1103 ( .A0(n4196), .A1(n4410), .B0(n1439), .B1(n4006), .Y(n1833) );
  AOI22X2 U1104 ( .A0(mem_rdata[26]), .A1(n4348), .B0(n4007), .B1(n1832), .Y(
        n1681) );
  OAI22XL U1105 ( .A0(n4196), .A1(n4411), .B0(n1434), .B1(n4006), .Y(n1832) );
  AOI22X2 U1106 ( .A0(mem_rdata[27]), .A1(n1345), .B0(n4007), .B1(n1831), .Y(
        n1680) );
  OAI22XL U1107 ( .A0(n4196), .A1(n4412), .B0(n1429), .B1(n4006), .Y(n1831) );
  AOI22X2 U1108 ( .A0(mem_rdata[28]), .A1(n1341), .B0(n4007), .B1(n1830), .Y(
        n1679) );
  OAI22XL U1109 ( .A0(n4195), .A1(n4413), .B0(n1424), .B1(n4006), .Y(n1830) );
  AOI22X2 U1110 ( .A0(mem_rdata[29]), .A1(n1345), .B0(n4007), .B1(n1829), .Y(
        n1678) );
  OAI22XL U1111 ( .A0(n4195), .A1(n4414), .B0(n1419), .B1(n4006), .Y(n1829) );
  AOI22X2 U1112 ( .A0(mem_rdata[30]), .A1(n1346), .B0(n4008), .B1(n1828), .Y(
        n1677) );
  OAI22XL U1113 ( .A0(n4195), .A1(n4416), .B0(n1409), .B1(n4006), .Y(n1828) );
  AOI22X2 U1114 ( .A0(mem_rdata[31]), .A1(n1348), .B0(n4008), .B1(n1827), .Y(
        n1676) );
  OAI22XL U1115 ( .A0(n4195), .A1(n4415), .B0(n1404), .B1(n4006), .Y(n1827) );
  AOI22X2 U1116 ( .A0(mem_rdata[32]), .A1(n1347), .B0(n4008), .B1(n1826), .Y(
        n1675) );
  OAI22XL U1117 ( .A0(n4197), .A1(n4417), .B0(n1522), .B1(n4003), .Y(n1826) );
  AOI22X2 U1118 ( .A0(mem_rdata[33]), .A1(n1343), .B0(n4008), .B1(n1825), .Y(
        n1674) );
  OAI22XL U1119 ( .A0(n4197), .A1(n4386), .B0(n1467), .B1(n4003), .Y(n1825) );
  AOI22X2 U1120 ( .A0(mem_rdata[34]), .A1(n1344), .B0(n4008), .B1(n1824), .Y(
        n1673) );
  OAI22XL U1121 ( .A0(n4197), .A1(n4387), .B0(n1412), .B1(n4003), .Y(n1824) );
  AOI22X2 U1122 ( .A0(mem_rdata[89]), .A1(n1346), .B0(n4012), .B1(n1767), .Y(
        n1618) );
  OAI22XL U1123 ( .A0(n4202), .A1(n4410), .B0(n1436), .B1(n1761), .Y(n1767) );
  AOI22X2 U1124 ( .A0(mem_rdata[90]), .A1(n1346), .B0(n4013), .B1(n1766), .Y(
        n1617) );
  OAI22XL U1125 ( .A0(n4203), .A1(n4411), .B0(n1431), .B1(n1761), .Y(n1766) );
  AOI22X2 U1126 ( .A0(mem_rdata[91]), .A1(n1346), .B0(n4014), .B1(n1765), .Y(
        n1616) );
  OAI22XL U1127 ( .A0(n4203), .A1(n4412), .B0(n1426), .B1(n1761), .Y(n1765) );
  AOI22X2 U1128 ( .A0(mem_rdata[92]), .A1(n1346), .B0(n4014), .B1(n1764), .Y(
        n1615) );
  OAI22XL U1129 ( .A0(n4203), .A1(n4413), .B0(n1421), .B1(n1761), .Y(n1764) );
  AOI22X2 U1130 ( .A0(mem_rdata[93]), .A1(n1346), .B0(n4014), .B1(n1763), .Y(
        n1614) );
  OAI22XL U1131 ( .A0(n4203), .A1(n4414), .B0(n1416), .B1(n1761), .Y(n1763) );
  AOI22X2 U1132 ( .A0(mem_rdata[94]), .A1(n1346), .B0(n4014), .B1(n1762), .Y(
        n1613) );
  OAI22XL U1133 ( .A0(n4203), .A1(n4416), .B0(n1406), .B1(n1761), .Y(n1762) );
  AOI22X2 U1134 ( .A0(mem_rdata[95]), .A1(n1346), .B0(n4014), .B1(n1760), .Y(
        n1612) );
  OAI22XL U1135 ( .A0(n4203), .A1(n4415), .B0(n1401), .B1(n1761), .Y(n1760) );
  AOI22X2 U1136 ( .A0(mem_rdata[96]), .A1(n1346), .B0(n4010), .B1(n1759), .Y(
        n1611) );
  OAI22XL U1137 ( .A0(n1525), .A1(n4005), .B0(n4191), .B1(n4417), .Y(n1759) );
  AOI22X2 U1138 ( .A0(mem_rdata[97]), .A1(n1346), .B0(n4008), .B1(n1758), .Y(
        n1610) );
  OAI22XL U1139 ( .A0(n1470), .A1(n4005), .B0(n4191), .B1(n4386), .Y(n1758) );
  AOI22X2 U1140 ( .A0(mem_rdata[98]), .A1(n1345), .B0(n4008), .B1(n1757), .Y(
        n1609) );
  OAI22XL U1141 ( .A0(n1415), .A1(n4005), .B0(n4191), .B1(n4387), .Y(n1757) );
  AOI22X2 U1142 ( .A0(mem_rdata[99]), .A1(n1345), .B0(n4007), .B1(n1756), .Y(
        n1608) );
  OAI22XL U1143 ( .A0(n1400), .A1(n4005), .B0(n4192), .B1(n4388), .Y(n1756) );
  AOI22X2 U1144 ( .A0(mem_rdata[100]), .A1(n1345), .B0(n4009), .B1(n1755), .Y(
        n1607) );
  OAI22XL U1145 ( .A0(n1395), .A1(n4005), .B0(n4192), .B1(n4389), .Y(n1755) );
  AOI22X2 U1146 ( .A0(mem_rdata[101]), .A1(n1345), .B0(n4011), .B1(n1754), .Y(
        n1606) );
  OAI22XL U1147 ( .A0(n1390), .A1(n4005), .B0(n4191), .B1(n4390), .Y(n1754) );
  AOI22X2 U1148 ( .A0(mem_rdata[102]), .A1(n1345), .B0(n4009), .B1(n1753), .Y(
        n1605) );
  OAI22XL U1149 ( .A0(n1385), .A1(n4005), .B0(n4191), .B1(n4391), .Y(n1753) );
  AOI22X2 U1150 ( .A0(mem_rdata[103]), .A1(n1345), .B0(n4014), .B1(n1752), .Y(
        n1604) );
  OAI22XL U1151 ( .A0(n1380), .A1(n4005), .B0(n4192), .B1(n4392), .Y(n1752) );
  AOI22X2 U1152 ( .A0(mem_rdata[104]), .A1(n1345), .B0(n4015), .B1(n1751), .Y(
        n1603) );
  OAI22XL U1153 ( .A0(n1375), .A1(n4005), .B0(n4192), .B1(n4393), .Y(n1751) );
  AOI22X2 U1154 ( .A0(mem_rdata[118]), .A1(n1344), .B0(n4013), .B1(n1737), .Y(
        n1589) );
  OAI22XL U1155 ( .A0(n1455), .A1(n4005), .B0(n4191), .B1(n4407), .Y(n1737) );
  AOI22X2 U1156 ( .A0(mem_rdata[119]), .A1(n1344), .B0(n4013), .B1(n1736), .Y(
        n1588) );
  OAI22XL U1157 ( .A0(n1450), .A1(n4005), .B0(n4193), .B1(n4408), .Y(n1736) );
  AOI22X2 U1158 ( .A0(mem_rdata[120]), .A1(n1344), .B0(n4013), .B1(n1735), .Y(
        n1587) );
  OAI22XL U1159 ( .A0(n1445), .A1(n1728), .B0(n4191), .B1(n4409), .Y(n1735) );
  AOI22X2 U1160 ( .A0(mem_rdata[121]), .A1(n1344), .B0(n4013), .B1(n1734), .Y(
        n1586) );
  OAI22XL U1161 ( .A0(n1440), .A1(n1728), .B0(n4193), .B1(n4410), .Y(n1734) );
  AOI22X2 U1162 ( .A0(mem_rdata[122]), .A1(n1343), .B0(n4013), .B1(n1733), .Y(
        n1585) );
  OAI22XL U1163 ( .A0(n1435), .A1(n1728), .B0(n4193), .B1(n4411), .Y(n1733) );
  AOI22X2 U1164 ( .A0(mem_rdata[123]), .A1(n1343), .B0(n4013), .B1(n1732), .Y(
        n1584) );
  OAI22XL U1165 ( .A0(n1430), .A1(n1728), .B0(n4193), .B1(n4412), .Y(n1732) );
  AOI22X2 U1166 ( .A0(mem_rdata[124]), .A1(n1343), .B0(n4013), .B1(n1731), .Y(
        n1583) );
  OAI22XL U1167 ( .A0(n1425), .A1(n1728), .B0(n4191), .B1(n4413), .Y(n1731) );
  AOI22X2 U1168 ( .A0(mem_rdata[125]), .A1(n1343), .B0(n4013), .B1(n1730), .Y(
        n1582) );
  OAI22XL U1169 ( .A0(n1420), .A1(n1728), .B0(n4193), .B1(n4414), .Y(n1730) );
  AOI22X2 U1170 ( .A0(mem_rdata[126]), .A1(n1343), .B0(n4015), .B1(n1729), .Y(
        n1581) );
  OAI22XL U1171 ( .A0(n1410), .A1(n1728), .B0(n4191), .B1(n4416), .Y(n1729) );
  AOI22X2 U1172 ( .A0(mem_rdata[127]), .A1(n1343), .B0(n4010), .B1(n1727), .Y(
        n1579) );
  OAI22XL U1173 ( .A0(n1405), .A1(n1728), .B0(n4193), .B1(n4415), .Y(n1727) );
  AOI22X2 U1174 ( .A0(mem_rdata[0]), .A1(n1343), .B0(n4012), .B1(n1726), .Y(
        n1545) );
  OAI22XL U1175 ( .A0(n4195), .A1(n4417), .B0(n1524), .B1(n1709), .Y(n1726) );
  AOI22X2 U1176 ( .A0(mem_rdata[1]), .A1(n1343), .B0(n4012), .B1(n1725), .Y(
        n1544) );
  OAI22XL U1177 ( .A0(n4195), .A1(n4386), .B0(n1469), .B1(n4006), .Y(n1725) );
  AOI22X2 U1178 ( .A0(mem_rdata[2]), .A1(n1343), .B0(n4008), .B1(n1724), .Y(
        n1543) );
  OAI22XL U1179 ( .A0(n4195), .A1(n4387), .B0(n1414), .B1(n4006), .Y(n1724) );
  AOI22X2 U1180 ( .A0(mem_rdata[3]), .A1(n1343), .B0(n4009), .B1(n1723), .Y(
        n1542) );
  OAI22XL U1181 ( .A0(n4195), .A1(n4388), .B0(n1399), .B1(n4006), .Y(n1723) );
  AOI22X2 U1182 ( .A0(mem_rdata[4]), .A1(n1343), .B0(n4015), .B1(n1722), .Y(
        n1541) );
  OAI22XL U1183 ( .A0(n4195), .A1(n4389), .B0(n1394), .B1(n4006), .Y(n1722) );
  AOI22X2 U1184 ( .A0(mem_rdata[5]), .A1(n1343), .B0(n1707), .B1(n1721), .Y(
        n1540) );
  OAI22XL U1185 ( .A0(n4195), .A1(n4390), .B0(n1389), .B1(n4006), .Y(n1721) );
  AOI22X2 U1186 ( .A0(mem_rdata[18]), .A1(n1349), .B0(n4007), .B1(n1840), .Y(
        n1689) );
  OAI22XL U1187 ( .A0(n4195), .A1(n4403), .B0(n1479), .B1(n4006), .Y(n1840) );
  AOI22X2 U1188 ( .A0(mem_rdata[35]), .A1(n1341), .B0(n4008), .B1(n1823), .Y(
        n1672) );
  OAI22XL U1189 ( .A0(n4197), .A1(n4388), .B0(n1397), .B1(n4003), .Y(n1823) );
  AOI22X2 U1190 ( .A0(mem_rdata[36]), .A1(n1348), .B0(n4008), .B1(n1822), .Y(
        n1671) );
  OAI22XL U1191 ( .A0(n4197), .A1(n4389), .B0(n1392), .B1(n4003), .Y(n1822) );
  AOI22X2 U1192 ( .A0(mem_rdata[37]), .A1(n1349), .B0(n4008), .B1(n1821), .Y(
        n1670) );
  OAI22XL U1193 ( .A0(n4197), .A1(n4390), .B0(n1387), .B1(n4003), .Y(n1821) );
  AOI22X2 U1194 ( .A0(mem_rdata[38]), .A1(n1342), .B0(n4008), .B1(n1820), .Y(
        n1669) );
  OAI22XL U1195 ( .A0(n10), .A1(n4391), .B0(n1382), .B1(n4003), .Y(n1820) );
  AOI22X2 U1196 ( .A0(mem_rdata[39]), .A1(n1342), .B0(n4008), .B1(n1819), .Y(
        n1668) );
  OAI22XL U1197 ( .A0(n10), .A1(n4392), .B0(n1377), .B1(n4003), .Y(n1819) );
  AOI22X2 U1198 ( .A0(mem_rdata[40]), .A1(n1342), .B0(n4008), .B1(n1818), .Y(
        n1667) );
  OAI22XL U1199 ( .A0(n10), .A1(n4393), .B0(n1372), .B1(n4003), .Y(n1818) );
  AOI22X2 U1200 ( .A0(mem_rdata[41]), .A1(n1342), .B0(n4008), .B1(n1817), .Y(
        n1666) );
  OAI22XL U1201 ( .A0(n10), .A1(n4394), .B0(n1364), .B1(n4003), .Y(n1817) );
  AOI22X2 U1202 ( .A0(mem_rdata[42]), .A1(n1342), .B0(n4009), .B1(n1816), .Y(
        n1665) );
  OAI22XL U1203 ( .A0(n10), .A1(n4395), .B0(n1517), .B1(n4003), .Y(n1816) );
  AOI22X2 U1204 ( .A0(mem_rdata[43]), .A1(n1342), .B0(n4009), .B1(n1815), .Y(
        n1664) );
  OAI22XL U1205 ( .A0(n10), .A1(n4396), .B0(n1512), .B1(n4003), .Y(n1815) );
  AOI22X2 U1206 ( .A0(mem_rdata[44]), .A1(n1342), .B0(n4009), .B1(n1814), .Y(
        n1663) );
  OAI22XL U1207 ( .A0(n4197), .A1(n4397), .B0(n1507), .B1(n1795), .Y(n1814) );
  AOI22X2 U1208 ( .A0(mem_rdata[45]), .A1(n1342), .B0(n4009), .B1(n1813), .Y(
        n1662) );
  OAI22XL U1209 ( .A0(n4197), .A1(n4398), .B0(n1502), .B1(n1795), .Y(n1813) );
  AOI22X2 U1210 ( .A0(mem_rdata[46]), .A1(n1342), .B0(n4009), .B1(n1812), .Y(
        n1661) );
  OAI22XL U1211 ( .A0(n4197), .A1(n4399), .B0(n1497), .B1(n1795), .Y(n1812) );
  AOI22X2 U1212 ( .A0(mem_rdata[47]), .A1(n1342), .B0(n4009), .B1(n1811), .Y(
        n1660) );
  OAI22XL U1213 ( .A0(n4197), .A1(n4400), .B0(n1492), .B1(n1795), .Y(n1811) );
  AOI22X2 U1214 ( .A0(mem_rdata[48]), .A1(n1342), .B0(n4009), .B1(n1810), .Y(
        n1659) );
  OAI22XL U1215 ( .A0(n4197), .A1(n4401), .B0(n1487), .B1(n1795), .Y(n1810) );
  AOI22X2 U1216 ( .A0(mem_rdata[49]), .A1(n1342), .B0(n4009), .B1(n1809), .Y(
        n1658) );
  OAI22XL U1217 ( .A0(n4198), .A1(n4402), .B0(n1482), .B1(n4003), .Y(n1809) );
  AOI22X2 U1218 ( .A0(mem_rdata[50]), .A1(n1348), .B0(n4009), .B1(n1808), .Y(
        n1657) );
  OAI22XL U1219 ( .A0(n4198), .A1(n4403), .B0(n1477), .B1(n4003), .Y(n1808) );
  AOI22X2 U1220 ( .A0(mem_rdata[51]), .A1(n1348), .B0(n4009), .B1(n1807), .Y(
        n1656) );
  OAI22XL U1221 ( .A0(n4198), .A1(n4404), .B0(n1472), .B1(n4003), .Y(n1807) );
  AOI22X2 U1222 ( .A0(mem_rdata[52]), .A1(n1348), .B0(n4009), .B1(n1806), .Y(
        n1655) );
  OAI22XL U1223 ( .A0(n4198), .A1(n4405), .B0(n1462), .B1(n4003), .Y(n1806) );
  AOI22X2 U1224 ( .A0(mem_rdata[53]), .A1(n1348), .B0(n4009), .B1(n1805), .Y(
        n1654) );
  OAI22XL U1225 ( .A0(n4198), .A1(n4406), .B0(n1457), .B1(n4003), .Y(n1805) );
  AOI22X2 U1226 ( .A0(mem_rdata[54]), .A1(n1348), .B0(n4010), .B1(n1804), .Y(
        n1653) );
  OAI22XL U1227 ( .A0(n4198), .A1(n4407), .B0(n1452), .B1(n4003), .Y(n1804) );
  AOI22X2 U1228 ( .A0(mem_rdata[55]), .A1(n1348), .B0(n4010), .B1(n1803), .Y(
        n1652) );
  OAI22XL U1229 ( .A0(n4198), .A1(n4408), .B0(n1447), .B1(n4003), .Y(n1803) );
  AOI22X2 U1230 ( .A0(mem_rdata[56]), .A1(n1348), .B0(n4010), .B1(n1802), .Y(
        n1651) );
  OAI22XL U1231 ( .A0(n4198), .A1(n4409), .B0(n1442), .B1(n1795), .Y(n1802) );
  AOI22X2 U1232 ( .A0(mem_rdata[57]), .A1(n1348), .B0(n4010), .B1(n1801), .Y(
        n1650) );
  OAI22XL U1233 ( .A0(n4198), .A1(n4410), .B0(n1437), .B1(n1795), .Y(n1801) );
  AOI22X2 U1234 ( .A0(mem_rdata[58]), .A1(n1348), .B0(n4010), .B1(n1800), .Y(
        n1649) );
  OAI22XL U1235 ( .A0(n4198), .A1(n4411), .B0(n1432), .B1(n1795), .Y(n1800) );
  AOI22X2 U1236 ( .A0(mem_rdata[59]), .A1(n1348), .B0(n4010), .B1(n1799), .Y(
        n1648) );
  OAI22XL U1237 ( .A0(n4198), .A1(n4412), .B0(n1427), .B1(n1795), .Y(n1799) );
  AOI22X2 U1238 ( .A0(mem_rdata[60]), .A1(n1348), .B0(n4010), .B1(n1798), .Y(
        n1647) );
  OAI22XL U1239 ( .A0(n4198), .A1(n4413), .B0(n1422), .B1(n1795), .Y(n1798) );
  AOI22X2 U1240 ( .A0(mem_rdata[61]), .A1(n1348), .B0(n4010), .B1(n1797), .Y(
        n1646) );
  OAI22XL U1241 ( .A0(n4198), .A1(n4414), .B0(n1417), .B1(n1795), .Y(n1797) );
  AOI22X2 U1242 ( .A0(mem_rdata[62]), .A1(n1347), .B0(n4010), .B1(n1796), .Y(
        n1645) );
  OAI22XL U1243 ( .A0(n4198), .A1(n4416), .B0(n1407), .B1(n1795), .Y(n1796) );
  AOI22X2 U1244 ( .A0(mem_rdata[63]), .A1(n1347), .B0(n4010), .B1(n1794), .Y(
        n1644) );
  OAI22XL U1245 ( .A0(n4198), .A1(n4415), .B0(n1402), .B1(n1795), .Y(n1794) );
  AOI22X2 U1246 ( .A0(mem_rdata[64]), .A1(n1347), .B0(n4010), .B1(n1792), .Y(
        n1643) );
  OAI22XL U1247 ( .A0(n4203), .A1(n4417), .B0(n1521), .B1(n4004), .Y(n1792) );
  AOI22X2 U1248 ( .A0(mem_rdata[65]), .A1(n1347), .B0(n4010), .B1(n1791), .Y(
        n1642) );
  OAI22XL U1249 ( .A0(n4203), .A1(n4386), .B0(n1466), .B1(n4004), .Y(n1791) );
  AOI22X2 U1250 ( .A0(mem_rdata[66]), .A1(n1347), .B0(n4011), .B1(n1790), .Y(
        n1641) );
  OAI22XL U1251 ( .A0(n4203), .A1(n4387), .B0(n1411), .B1(n4004), .Y(n1790) );
  AOI22X2 U1252 ( .A0(mem_rdata[67]), .A1(n1347), .B0(n4011), .B1(n1789), .Y(
        n1640) );
  OAI22XL U1253 ( .A0(n4203), .A1(n4388), .B0(n1396), .B1(n4004), .Y(n1789) );
  AOI22X2 U1254 ( .A0(mem_rdata[68]), .A1(n1347), .B0(n4011), .B1(n1788), .Y(
        n1639) );
  OAI22XL U1255 ( .A0(n4203), .A1(n4389), .B0(n1391), .B1(n4004), .Y(n1788) );
  AOI22X2 U1256 ( .A0(mem_rdata[69]), .A1(n1347), .B0(n4011), .B1(n1787), .Y(
        n1638) );
  OAI22XL U1257 ( .A0(n4203), .A1(n4390), .B0(n1386), .B1(n4004), .Y(n1787) );
  AOI22X2 U1258 ( .A0(mem_rdata[70]), .A1(n1347), .B0(n4011), .B1(n1786), .Y(
        n1637) );
  OAI22XL U1259 ( .A0(n4202), .A1(n4391), .B0(n1381), .B1(n4004), .Y(n1786) );
  AOI22X2 U1260 ( .A0(mem_rdata[71]), .A1(n1347), .B0(n4011), .B1(n1785), .Y(
        n1636) );
  OAI22XL U1261 ( .A0(n4203), .A1(n4392), .B0(n1376), .B1(n4004), .Y(n1785) );
  AOI22X2 U1262 ( .A0(mem_rdata[72]), .A1(n1347), .B0(n4011), .B1(n1784), .Y(
        n1635) );
  OAI22XL U1263 ( .A0(n4203), .A1(n4393), .B0(n1371), .B1(n4004), .Y(n1784) );
  AOI22X2 U1264 ( .A0(mem_rdata[73]), .A1(n1347), .B0(n4011), .B1(n1783), .Y(
        n1634) );
  OAI22XL U1265 ( .A0(n4202), .A1(n4394), .B0(n1362), .B1(n4004), .Y(n1783) );
  AOI22X2 U1266 ( .A0(mem_rdata[74]), .A1(n1347), .B0(n4011), .B1(n1782), .Y(
        n1633) );
  OAI22XL U1267 ( .A0(n4202), .A1(n4395), .B0(n1516), .B1(n4004), .Y(n1782) );
  AOI22X2 U1268 ( .A0(mem_rdata[75]), .A1(n1346), .B0(n4011), .B1(n1781), .Y(
        n1632) );
  OAI22XL U1269 ( .A0(n4202), .A1(n4396), .B0(n1511), .B1(n4004), .Y(n1781) );
  AOI22X2 U1270 ( .A0(mem_rdata[76]), .A1(n1348), .B0(n4011), .B1(n1780), .Y(
        n1631) );
  OAI22XL U1271 ( .A0(n4202), .A1(n4397), .B0(n1506), .B1(n1761), .Y(n1780) );
  AOI22X2 U1272 ( .A0(mem_rdata[77]), .A1(n1347), .B0(n4011), .B1(n1779), .Y(
        n1630) );
  OAI22XL U1273 ( .A0(n4202), .A1(n4398), .B0(n1501), .B1(n1761), .Y(n1779) );
  AOI22X2 U1274 ( .A0(mem_rdata[78]), .A1(n1346), .B0(n4012), .B1(n1778), .Y(
        n1629) );
  OAI22XL U1275 ( .A0(n4202), .A1(n4399), .B0(n1496), .B1(n1761), .Y(n1778) );
  AOI22X2 U1276 ( .A0(mem_rdata[79]), .A1(n1345), .B0(n4012), .B1(n1777), .Y(
        n1628) );
  OAI22XL U1277 ( .A0(n4202), .A1(n4400), .B0(n1491), .B1(n1761), .Y(n1777) );
  AOI22X2 U1278 ( .A0(mem_rdata[80]), .A1(n1349), .B0(n4012), .B1(n1776), .Y(
        n1627) );
  OAI22XL U1279 ( .A0(n4202), .A1(n4401), .B0(n1486), .B1(n1761), .Y(n1776) );
  AOI22X2 U1280 ( .A0(mem_rdata[81]), .A1(n1342), .B0(n4012), .B1(n1775), .Y(
        n1626) );
  OAI22XL U1281 ( .A0(n4202), .A1(n4402), .B0(n1481), .B1(n4004), .Y(n1775) );
  AOI22X2 U1282 ( .A0(mem_rdata[82]), .A1(n1342), .B0(n4012), .B1(n1774), .Y(
        n1625) );
  OAI22XL U1283 ( .A0(n4202), .A1(n4403), .B0(n1476), .B1(n4004), .Y(n1774) );
  AOI22X2 U1284 ( .A0(mem_rdata[83]), .A1(n4348), .B0(n4012), .B1(n1773), .Y(
        n1624) );
  OAI22XL U1285 ( .A0(n4202), .A1(n4404), .B0(n1471), .B1(n4004), .Y(n1773) );
  AOI22X2 U1286 ( .A0(mem_rdata[84]), .A1(n4348), .B0(n4012), .B1(n1772), .Y(
        n1623) );
  OAI22XL U1287 ( .A0(n4202), .A1(n4405), .B0(n1461), .B1(n4004), .Y(n1772) );
  AOI22X2 U1288 ( .A0(mem_rdata[85]), .A1(n4348), .B0(n4012), .B1(n1771), .Y(
        n1622) );
  OAI22XL U1289 ( .A0(n4202), .A1(n4406), .B0(n1456), .B1(n4004), .Y(n1771) );
  AOI22X2 U1290 ( .A0(mem_rdata[86]), .A1(n1346), .B0(n4012), .B1(n1770), .Y(
        n1621) );
  OAI22XL U1291 ( .A0(n4202), .A1(n4407), .B0(n1451), .B1(n4004), .Y(n1770) );
  AOI22X2 U1292 ( .A0(mem_rdata[87]), .A1(n1346), .B0(n4012), .B1(n1769), .Y(
        n1620) );
  OAI22XL U1293 ( .A0(n4202), .A1(n4408), .B0(n1446), .B1(n4004), .Y(n1769) );
  AOI22X2 U1294 ( .A0(mem_rdata[88]), .A1(n1346), .B0(n4012), .B1(n1768), .Y(
        n1619) );
  OAI22XL U1295 ( .A0(n4202), .A1(n4409), .B0(n1441), .B1(n1761), .Y(n1768) );
  AOI22X2 U1296 ( .A0(mem_rdata[105]), .A1(n1345), .B0(n4007), .B1(n1750), .Y(
        n1602) );
  OAI22XL U1297 ( .A0(n1369), .A1(n4005), .B0(n4192), .B1(n4394), .Y(n1750) );
  AOI22X2 U1298 ( .A0(mem_rdata[106]), .A1(n1345), .B0(n4014), .B1(n1749), .Y(
        n1601) );
  OAI22XL U1299 ( .A0(n1520), .A1(n4005), .B0(n4192), .B1(n4395), .Y(n1749) );
  AOI22X2 U1300 ( .A0(mem_rdata[107]), .A1(n1345), .B0(n4007), .B1(n1748), .Y(
        n1600) );
  OAI22XL U1301 ( .A0(n1515), .A1(n4005), .B0(n4192), .B1(n4396), .Y(n1748) );
  AOI22X2 U1302 ( .A0(mem_rdata[108]), .A1(n1345), .B0(n4013), .B1(n1747), .Y(
        n1599) );
  OAI22XL U1303 ( .A0(n1510), .A1(n1728), .B0(n4192), .B1(n4397), .Y(n1747) );
  AOI22X2 U1304 ( .A0(mem_rdata[109]), .A1(n1345), .B0(n4010), .B1(n1746), .Y(
        n1598) );
  OAI22XL U1305 ( .A0(n1505), .A1(n1728), .B0(n4192), .B1(n4398), .Y(n1746) );
  AOI22X2 U1306 ( .A0(mem_rdata[110]), .A1(n1344), .B0(n4015), .B1(n1745), .Y(
        n1597) );
  OAI22XL U1307 ( .A0(n1500), .A1(n1728), .B0(n4192), .B1(n4399), .Y(n1745) );
  AOI22X2 U1308 ( .A0(mem_rdata[111]), .A1(n1344), .B0(n4015), .B1(n1744), .Y(
        n1596) );
  OAI22XL U1309 ( .A0(n1495), .A1(n1728), .B0(n4192), .B1(n4400), .Y(n1744) );
  AOI22X2 U1310 ( .A0(mem_rdata[112]), .A1(n1344), .B0(n4015), .B1(n1743), .Y(
        n1595) );
  OAI22XL U1311 ( .A0(n1490), .A1(n1728), .B0(n4192), .B1(n4401), .Y(n1743) );
  AOI22X2 U1312 ( .A0(mem_rdata[113]), .A1(n1344), .B0(n1707), .B1(n1742), .Y(
        n1594) );
  OAI22XL U1313 ( .A0(n1485), .A1(n4005), .B0(n4192), .B1(n4402), .Y(n1742) );
  AOI22X2 U1314 ( .A0(mem_rdata[114]), .A1(n1344), .B0(n4013), .B1(n1741), .Y(
        n1593) );
  OAI22XL U1315 ( .A0(n1480), .A1(n4005), .B0(n4192), .B1(n4403), .Y(n1741) );
  AOI22X2 U1316 ( .A0(mem_rdata[115]), .A1(n1344), .B0(n4013), .B1(n1740), .Y(
        n1592) );
  OAI22XL U1317 ( .A0(n1475), .A1(n4005), .B0(n4192), .B1(n4404), .Y(n1740) );
  AOI22X2 U1318 ( .A0(mem_rdata[116]), .A1(n1344), .B0(n4013), .B1(n1739), .Y(
        n1591) );
  OAI22XL U1319 ( .A0(n1465), .A1(n4005), .B0(n4193), .B1(n4405), .Y(n1739) );
  AOI22X2 U1320 ( .A0(mem_rdata[117]), .A1(n1344), .B0(n4013), .B1(n1738), .Y(
        n1590) );
  OAI22XL U1321 ( .A0(n1460), .A1(n4005), .B0(n4191), .B1(n4406), .Y(n1738) );
  AOI22X2 U1322 ( .A0(mem_rdata[6]), .A1(n1341), .B0(n4013), .B1(n1720), .Y(
        n1539) );
  OAI22XL U1323 ( .A0(n4194), .A1(n4391), .B0(n1384), .B1(n1709), .Y(n1720) );
  AOI22X2 U1324 ( .A0(mem_rdata[7]), .A1(n1341), .B0(n4011), .B1(n1719), .Y(
        n1538) );
  OAI22XL U1325 ( .A0(n4194), .A1(n4392), .B0(n1379), .B1(n1709), .Y(n1719) );
  AOI22X2 U1326 ( .A0(mem_rdata[8]), .A1(n1341), .B0(n4015), .B1(n1718), .Y(
        n1537) );
  OAI22XL U1327 ( .A0(n4194), .A1(n4393), .B0(n1374), .B1(n1709), .Y(n1718) );
  AOI22X2 U1328 ( .A0(mem_rdata[9]), .A1(n1341), .B0(n4015), .B1(n1717), .Y(
        n1536) );
  OAI22XL U1329 ( .A0(n4194), .A1(n4394), .B0(n1367), .B1(n1709), .Y(n1717) );
  AOI22X2 U1330 ( .A0(mem_rdata[10]), .A1(n1341), .B0(n4014), .B1(n1716), .Y(
        n1535) );
  OAI22XL U1331 ( .A0(n4194), .A1(n4395), .B0(n1519), .B1(n1709), .Y(n1716) );
  AOI22X2 U1332 ( .A0(mem_rdata[11]), .A1(n1341), .B0(n4014), .B1(n1715), .Y(
        n1534) );
  OAI22XL U1333 ( .A0(n4194), .A1(n4396), .B0(n1514), .B1(n1709), .Y(n1715) );
  AOI22X2 U1334 ( .A0(mem_rdata[12]), .A1(n1341), .B0(n4014), .B1(n1714), .Y(
        n1533) );
  OAI22XL U1335 ( .A0(n4194), .A1(n4397), .B0(n1509), .B1(n1709), .Y(n1714) );
  AOI22X2 U1336 ( .A0(mem_rdata[13]), .A1(n1341), .B0(n4014), .B1(n1713), .Y(
        n1532) );
  OAI22XL U1337 ( .A0(n4194), .A1(n4398), .B0(n1504), .B1(n1709), .Y(n1713) );
  AOI22X2 U1338 ( .A0(mem_rdata[14]), .A1(n1341), .B0(n4014), .B1(n1712), .Y(
        n1531) );
  OAI22XL U1339 ( .A0(n4194), .A1(n4399), .B0(n1499), .B1(n1709), .Y(n1712) );
  AOI22X2 U1340 ( .A0(mem_rdata[15]), .A1(n1341), .B0(n4014), .B1(n1711), .Y(
        n1530) );
  OAI22XL U1341 ( .A0(n4194), .A1(n4400), .B0(n1494), .B1(n1709), .Y(n1711) );
  AOI22X2 U1342 ( .A0(mem_rdata[16]), .A1(n1341), .B0(n4014), .B1(n1710), .Y(
        n1529) );
  OAI22XL U1343 ( .A0(n4194), .A1(n4401), .B0(n1489), .B1(n1709), .Y(n1710) );
  AOI22X2 U1344 ( .A0(mem_rdata[17]), .A1(n1341), .B0(n4014), .B1(n1708), .Y(
        n1527) );
  OAI22XL U1345 ( .A0(n4194), .A1(n4402), .B0(n1484), .B1(n1709), .Y(n1708) );
  XOR2XL U1346 ( .A(\tag_r[1][3] ), .B(proc_addr[8]), .Y(n2034) );
  XOR2XL U1347 ( .A(\tag_r[1][17] ), .B(proc_addr[22]), .Y(n2042) );
  XOR2XL U1348 ( .A(\tag_r[2][3] ), .B(proc_addr[8]), .Y(n2067) );
  XOR2XL U1349 ( .A(\tag_r[2][17] ), .B(proc_addr[22]), .Y(n2075) );
  XOR2XL U1350 ( .A(\tag_r[3][3] ), .B(proc_addr[8]), .Y(n2100) );
  XOR2XL U1351 ( .A(\tag_r[3][17] ), .B(proc_addr[22]), .Y(n2108) );
  XOR2XL U1352 ( .A(\tag_r[0][3] ), .B(proc_addr[8]), .Y(n2001) );
  XOR2XL U1353 ( .A(\tag_r[0][17] ), .B(proc_addr[22]), .Y(n2009) );
  XOR2XL U1354 ( .A(\tag_r[5][3] ), .B(proc_addr[8]), .Y(n1898) );
  XOR2XL U1355 ( .A(\tag_r[5][17] ), .B(proc_addr[22]), .Y(n1906) );
  XOR2XL U1356 ( .A(\tag_r[6][3] ), .B(proc_addr[8]), .Y(n1931) );
  XOR2XL U1357 ( .A(\tag_r[6][17] ), .B(proc_addr[22]), .Y(n1939) );
  XOR2XL U1358 ( .A(\tag_r[7][3] ), .B(proc_addr[8]), .Y(n1964) );
  XOR2XL U1359 ( .A(\tag_r[7][17] ), .B(proc_addr[22]), .Y(n1972) );
  XOR2XL U1360 ( .A(\tag_r[4][3] ), .B(proc_addr[8]), .Y(n1865) );
  XOR2XL U1361 ( .A(\tag_r[4][17] ), .B(proc_addr[22]), .Y(n1873) );
  NOR3X1 U1362 ( .A(n2024), .B(n2025), .C(n2026), .Y(n2023) );
  XOR2XL U1363 ( .A(\tag_r[1][14] ), .B(proc_addr[19]), .Y(n2026) );
  XOR2XL U1364 ( .A(\tag_r[1][15] ), .B(proc_addr[20]), .Y(n2024) );
  XOR2XL U1365 ( .A(\tag_r[1][13] ), .B(proc_addr[18]), .Y(n2025) );
  NOR3X1 U1366 ( .A(n2057), .B(n2058), .C(n2059), .Y(n2056) );
  XOR2XL U1367 ( .A(\tag_r[2][14] ), .B(proc_addr[19]), .Y(n2059) );
  XOR2XL U1368 ( .A(\tag_r[2][15] ), .B(proc_addr[20]), .Y(n2057) );
  XOR2XL U1369 ( .A(\tag_r[2][13] ), .B(proc_addr[18]), .Y(n2058) );
  NOR3X1 U1370 ( .A(n2090), .B(n2091), .C(n2092), .Y(n2089) );
  XOR2XL U1371 ( .A(\tag_r[3][14] ), .B(proc_addr[19]), .Y(n2092) );
  XOR2XL U1372 ( .A(\tag_r[3][15] ), .B(proc_addr[20]), .Y(n2090) );
  XOR2XL U1373 ( .A(\tag_r[3][13] ), .B(proc_addr[18]), .Y(n2091) );
  NOR3X1 U1374 ( .A(n1991), .B(n1992), .C(n1993), .Y(n1990) );
  XOR2XL U1375 ( .A(\tag_r[0][14] ), .B(proc_addr[19]), .Y(n1993) );
  XOR2XL U1376 ( .A(\tag_r[0][15] ), .B(proc_addr[20]), .Y(n1991) );
  XOR2XL U1377 ( .A(\tag_r[0][13] ), .B(proc_addr[18]), .Y(n1992) );
  NOR3X1 U1378 ( .A(n1888), .B(n1889), .C(n1890), .Y(n1887) );
  XOR2XL U1379 ( .A(\tag_r[5][14] ), .B(proc_addr[19]), .Y(n1890) );
  XOR2XL U1380 ( .A(\tag_r[5][15] ), .B(proc_addr[20]), .Y(n1888) );
  XOR2XL U1381 ( .A(\tag_r[5][13] ), .B(proc_addr[18]), .Y(n1889) );
  NOR3X1 U1382 ( .A(n1921), .B(n1922), .C(n1923), .Y(n1920) );
  XOR2XL U1383 ( .A(\tag_r[6][14] ), .B(proc_addr[19]), .Y(n1923) );
  XOR2XL U1384 ( .A(\tag_r[6][15] ), .B(proc_addr[20]), .Y(n1921) );
  XOR2XL U1385 ( .A(\tag_r[6][13] ), .B(proc_addr[18]), .Y(n1922) );
  NOR3X1 U1386 ( .A(n1954), .B(n1955), .C(n1956), .Y(n1953) );
  XOR2XL U1387 ( .A(\tag_r[7][14] ), .B(proc_addr[19]), .Y(n1956) );
  XOR2XL U1388 ( .A(\tag_r[7][15] ), .B(proc_addr[20]), .Y(n1954) );
  XOR2XL U1389 ( .A(\tag_r[7][13] ), .B(proc_addr[18]), .Y(n1955) );
  NOR3X1 U1390 ( .A(n1855), .B(n1856), .C(n1857), .Y(n1854) );
  XOR2XL U1391 ( .A(\tag_r[4][14] ), .B(proc_addr[19]), .Y(n1857) );
  XOR2XL U1392 ( .A(\tag_r[4][15] ), .B(proc_addr[20]), .Y(n1855) );
  XOR2XL U1393 ( .A(\tag_r[4][13] ), .B(proc_addr[18]), .Y(n1856) );
  XOR2XL U1394 ( .A(n1254), .B(proc_addr[14]), .Y(n2029) );
  XOR2XL U1395 ( .A(n1240), .B(proc_addr[28]), .Y(n2037) );
  XOR2XL U1396 ( .A(n1242), .B(proc_addr[26]), .Y(n2022) );
  XOR2XL U1397 ( .A(n1229), .B(proc_addr[14]), .Y(n2062) );
  XOR2XL U1398 ( .A(n1215), .B(proc_addr[28]), .Y(n2070) );
  XOR2XL U1399 ( .A(n1217), .B(proc_addr[26]), .Y(n2055) );
  XOR2XL U1400 ( .A(n1204), .B(proc_addr[14]), .Y(n2095) );
  XOR2XL U1401 ( .A(n1190), .B(proc_addr[28]), .Y(n2103) );
  XOR2XL U1402 ( .A(n1192), .B(proc_addr[26]), .Y(n2088) );
  XOR2XL U1403 ( .A(n1265), .B(proc_addr[28]), .Y(n2004) );
  XOR2XL U1404 ( .A(n1267), .B(proc_addr[26]), .Y(n1989) );
  XOR2XL U1405 ( .A(n1272), .B(proc_addr[21]), .Y(n2012) );
  XOR2XL U1406 ( .A(n1154), .B(proc_addr[14]), .Y(n1893) );
  XOR2XL U1407 ( .A(n1140), .B(proc_addr[28]), .Y(n1901) );
  XOR2XL U1408 ( .A(n1142), .B(proc_addr[26]), .Y(n1886) );
  XOR2XL U1409 ( .A(n1129), .B(proc_addr[14]), .Y(n1926) );
  XOR2XL U1410 ( .A(n1115), .B(proc_addr[28]), .Y(n1934) );
  XOR2XL U1411 ( .A(n1117), .B(proc_addr[26]), .Y(n1919) );
  XOR2XL U1412 ( .A(n1104), .B(proc_addr[14]), .Y(n1959) );
  XOR2XL U1413 ( .A(n1090), .B(proc_addr[28]), .Y(n1967) );
  XOR2XL U1414 ( .A(n1092), .B(proc_addr[26]), .Y(n1952) );
  XOR2XL U1415 ( .A(n1256), .B(proc_addr[12]), .Y(n2028) );
  XOR2XL U1416 ( .A(n1241), .B(proc_addr[27]), .Y(n2036) );
  XOR2XL U1417 ( .A(n1244), .B(proc_addr[24]), .Y(n2021) );
  XOR2XL U1418 ( .A(n1231), .B(proc_addr[12]), .Y(n2061) );
  XOR2XL U1419 ( .A(n1216), .B(proc_addr[27]), .Y(n2069) );
  XOR2XL U1420 ( .A(n1219), .B(proc_addr[24]), .Y(n2054) );
  XOR2XL U1421 ( .A(n1206), .B(proc_addr[12]), .Y(n2094) );
  XOR2XL U1422 ( .A(n1191), .B(proc_addr[27]), .Y(n2102) );
  XOR2XL U1423 ( .A(n1194), .B(proc_addr[24]), .Y(n2087) );
  XOR2XL U1424 ( .A(n1266), .B(proc_addr[27]), .Y(n2003) );
  XOR2XL U1425 ( .A(n1269), .B(proc_addr[24]), .Y(n1988) );
  XOR2XL U1426 ( .A(n1283), .B(proc_addr[10]), .Y(n2011) );
  XOR2XL U1427 ( .A(n1156), .B(proc_addr[12]), .Y(n1892) );
  XOR2XL U1428 ( .A(n1141), .B(proc_addr[27]), .Y(n1900) );
  XOR2XL U1429 ( .A(n1144), .B(proc_addr[24]), .Y(n1885) );
  XOR2XL U1430 ( .A(n1131), .B(proc_addr[12]), .Y(n1925) );
  XOR2XL U1431 ( .A(n1116), .B(proc_addr[27]), .Y(n1933) );
  XOR2XL U1432 ( .A(n1119), .B(proc_addr[24]), .Y(n1918) );
  XOR2XL U1433 ( .A(n1106), .B(proc_addr[12]), .Y(n1958) );
  XOR2XL U1434 ( .A(n1091), .B(proc_addr[27]), .Y(n1966) );
  XOR2XL U1435 ( .A(n1094), .B(proc_addr[24]), .Y(n1951) );
  XOR2XL U1436 ( .A(n1255), .B(proc_addr[13]), .Y(n2027) );
  XOR2XL U1437 ( .A(n1239), .B(proc_addr[29]), .Y(n2035) );
  XOR2XL U1438 ( .A(n1243), .B(proc_addr[25]), .Y(n2020) );
  XOR2XL U1439 ( .A(n1230), .B(proc_addr[13]), .Y(n2060) );
  XOR2XL U1440 ( .A(n1214), .B(proc_addr[29]), .Y(n2068) );
  XOR2XL U1441 ( .A(n1218), .B(proc_addr[25]), .Y(n2053) );
  XOR2XL U1442 ( .A(n1205), .B(proc_addr[13]), .Y(n2093) );
  XOR2XL U1443 ( .A(n1189), .B(proc_addr[29]), .Y(n2101) );
  XOR2XL U1444 ( .A(n1193), .B(proc_addr[25]), .Y(n2086) );
  XOR2XL U1445 ( .A(n1264), .B(proc_addr[29]), .Y(n2002) );
  XOR2XL U1446 ( .A(n1268), .B(proc_addr[25]), .Y(n1987) );
  XOR2XL U1447 ( .A(n1278), .B(proc_addr[15]), .Y(n2010) );
  XOR2XL U1448 ( .A(n1155), .B(proc_addr[13]), .Y(n1891) );
  XOR2XL U1449 ( .A(n1139), .B(proc_addr[29]), .Y(n1899) );
  XOR2XL U1450 ( .A(n1143), .B(proc_addr[25]), .Y(n1884) );
  XOR2XL U1451 ( .A(n1130), .B(proc_addr[13]), .Y(n1924) );
  XOR2XL U1452 ( .A(n1114), .B(proc_addr[29]), .Y(n1932) );
  XOR2XL U1453 ( .A(n1118), .B(proc_addr[25]), .Y(n1917) );
  XOR2XL U1454 ( .A(n1105), .B(proc_addr[13]), .Y(n1957) );
  XOR2XL U1455 ( .A(n1089), .B(proc_addr[29]), .Y(n1965) );
  XOR2XL U1456 ( .A(n1093), .B(proc_addr[25]), .Y(n1950) );
  NOR4X1 U1457 ( .A(n2031), .B(n2032), .C(n2033), .D(n2034), .Y(n2030) );
  XOR2XL U1458 ( .A(\tag_r[1][0] ), .B(proc_addr[5]), .Y(n2031) );
  XOR2XL U1459 ( .A(\tag_r[1][1] ), .B(proc_addr[6]), .Y(n2032) );
  XOR2XL U1460 ( .A(\tag_r[1][2] ), .B(proc_addr[7]), .Y(n2033) );
  NOR4X1 U1461 ( .A(n2039), .B(n2040), .C(n2041), .D(n2042), .Y(n2038) );
  XOR2XL U1462 ( .A(\tag_r[1][12] ), .B(proc_addr[17]), .Y(n2039) );
  XOR2XL U1463 ( .A(\tag_r[1][16] ), .B(proc_addr[21]), .Y(n2040) );
  XOR2XL U1464 ( .A(\tag_r[1][18] ), .B(proc_addr[23]), .Y(n2041) );
  NOR4X1 U1465 ( .A(n2064), .B(n2065), .C(n2066), .D(n2067), .Y(n2063) );
  XOR2XL U1466 ( .A(\tag_r[2][0] ), .B(proc_addr[5]), .Y(n2064) );
  XOR2XL U1467 ( .A(\tag_r[2][1] ), .B(proc_addr[6]), .Y(n2065) );
  XOR2XL U1468 ( .A(\tag_r[2][2] ), .B(proc_addr[7]), .Y(n2066) );
  NOR4X1 U1469 ( .A(n2072), .B(n2073), .C(n2074), .D(n2075), .Y(n2071) );
  XOR2XL U1470 ( .A(\tag_r[2][12] ), .B(proc_addr[17]), .Y(n2072) );
  XOR2XL U1471 ( .A(\tag_r[2][16] ), .B(proc_addr[21]), .Y(n2073) );
  XOR2XL U1472 ( .A(\tag_r[2][18] ), .B(proc_addr[23]), .Y(n2074) );
  NOR4X1 U1473 ( .A(n2097), .B(n2098), .C(n2099), .D(n2100), .Y(n2096) );
  XOR2XL U1474 ( .A(\tag_r[3][0] ), .B(proc_addr[5]), .Y(n2097) );
  XOR2XL U1475 ( .A(\tag_r[3][1] ), .B(proc_addr[6]), .Y(n2098) );
  XOR2XL U1476 ( .A(\tag_r[3][2] ), .B(proc_addr[7]), .Y(n2099) );
  NOR4X1 U1477 ( .A(n2105), .B(n2106), .C(n2107), .D(n2108), .Y(n2104) );
  XOR2XL U1478 ( .A(\tag_r[3][12] ), .B(proc_addr[17]), .Y(n2105) );
  XOR2XL U1479 ( .A(\tag_r[3][16] ), .B(proc_addr[21]), .Y(n2106) );
  XOR2XL U1480 ( .A(\tag_r[3][18] ), .B(proc_addr[23]), .Y(n2107) );
  NOR4X1 U1481 ( .A(n1998), .B(n1999), .C(n2000), .D(n2001), .Y(n1997) );
  XOR2XL U1482 ( .A(\tag_r[0][0] ), .B(proc_addr[5]), .Y(n1998) );
  XOR2XL U1483 ( .A(\tag_r[0][1] ), .B(proc_addr[6]), .Y(n1999) );
  XOR2XL U1484 ( .A(\tag_r[0][2] ), .B(proc_addr[7]), .Y(n2000) );
  NOR4X1 U1485 ( .A(n2006), .B(n2007), .C(n2008), .D(n2009), .Y(n2005) );
  XOR2XL U1486 ( .A(\tag_r[0][12] ), .B(proc_addr[17]), .Y(n2006) );
  XOR2XL U1487 ( .A(\tag_r[0][11] ), .B(proc_addr[16]), .Y(n2007) );
  XOR2XL U1488 ( .A(\tag_r[0][18] ), .B(proc_addr[23]), .Y(n2008) );
  NOR4X1 U1489 ( .A(n1895), .B(n1896), .C(n1897), .D(n1898), .Y(n1894) );
  XOR2XL U1490 ( .A(\tag_r[5][0] ), .B(proc_addr[5]), .Y(n1895) );
  XOR2XL U1491 ( .A(\tag_r[5][1] ), .B(proc_addr[6]), .Y(n1896) );
  XOR2XL U1492 ( .A(\tag_r[5][2] ), .B(proc_addr[7]), .Y(n1897) );
  NOR4X1 U1493 ( .A(n1903), .B(n1904), .C(n1905), .D(n1906), .Y(n1902) );
  XOR2XL U1494 ( .A(\tag_r[5][12] ), .B(proc_addr[17]), .Y(n1903) );
  XOR2XL U1495 ( .A(\tag_r[5][16] ), .B(proc_addr[21]), .Y(n1904) );
  XOR2XL U1496 ( .A(\tag_r[5][18] ), .B(proc_addr[23]), .Y(n1905) );
  NOR4X1 U1497 ( .A(n1928), .B(n1929), .C(n1930), .D(n1931), .Y(n1927) );
  XOR2XL U1498 ( .A(\tag_r[6][0] ), .B(proc_addr[5]), .Y(n1928) );
  XOR2XL U1499 ( .A(\tag_r[6][1] ), .B(proc_addr[6]), .Y(n1929) );
  XOR2XL U1500 ( .A(\tag_r[6][2] ), .B(proc_addr[7]), .Y(n1930) );
  NOR4X1 U1501 ( .A(n1936), .B(n1937), .C(n1938), .D(n1939), .Y(n1935) );
  XOR2XL U1502 ( .A(\tag_r[6][12] ), .B(proc_addr[17]), .Y(n1936) );
  XOR2XL U1503 ( .A(\tag_r[6][16] ), .B(proc_addr[21]), .Y(n1937) );
  XOR2XL U1504 ( .A(\tag_r[6][18] ), .B(proc_addr[23]), .Y(n1938) );
  NOR4X1 U1505 ( .A(n1961), .B(n1962), .C(n1963), .D(n1964), .Y(n1960) );
  XOR2XL U1506 ( .A(\tag_r[7][0] ), .B(proc_addr[5]), .Y(n1961) );
  XOR2XL U1507 ( .A(\tag_r[7][1] ), .B(proc_addr[6]), .Y(n1962) );
  XOR2XL U1508 ( .A(\tag_r[7][2] ), .B(proc_addr[7]), .Y(n1963) );
  NOR4X1 U1509 ( .A(n1969), .B(n1970), .C(n1971), .D(n1972), .Y(n1968) );
  XOR2XL U1510 ( .A(\tag_r[7][12] ), .B(proc_addr[17]), .Y(n1969) );
  XOR2XL U1511 ( .A(\tag_r[7][11] ), .B(proc_addr[16]), .Y(n1970) );
  XOR2XL U1512 ( .A(\tag_r[7][18] ), .B(proc_addr[23]), .Y(n1971) );
  NOR4X1 U1513 ( .A(n1862), .B(n1863), .C(n1864), .D(n1865), .Y(n1861) );
  XOR2XL U1514 ( .A(\tag_r[4][0] ), .B(proc_addr[5]), .Y(n1862) );
  XOR2XL U1515 ( .A(\tag_r[4][1] ), .B(proc_addr[6]), .Y(n1863) );
  XOR2XL U1516 ( .A(\tag_r[4][2] ), .B(proc_addr[7]), .Y(n1864) );
  NOR4X1 U1517 ( .A(n1870), .B(n1871), .C(n1872), .D(n1873), .Y(n1869) );
  XOR2XL U1518 ( .A(\tag_r[4][12] ), .B(proc_addr[17]), .Y(n1870) );
  XOR2XL U1519 ( .A(\tag_r[4][16] ), .B(proc_addr[21]), .Y(n1871) );
  XOR2XL U1520 ( .A(\tag_r[4][18] ), .B(proc_addr[23]), .Y(n1872) );
  NOR4X1 U1521 ( .A(n2628), .B(n50), .C(n2014), .D(n2015), .Y(n2013) );
  XOR2XL U1522 ( .A(\tag_r[0][4] ), .B(proc_addr[9]), .Y(n2014) );
  XOR2XL U1523 ( .A(\tag_r[0][6] ), .B(proc_addr[11]), .Y(n2015) );
  NOR4X1 U1524 ( .A(n4141), .B(n43), .C(n1977), .D(n1978), .Y(n1976) );
  XOR2XL U1525 ( .A(\tag_r[7][4] ), .B(proc_addr[9]), .Y(n1977) );
  XOR2XL U1526 ( .A(\tag_r[7][6] ), .B(proc_addr[11]), .Y(n1978) );
  NOR4X1 U1527 ( .A(n4112), .B(n46), .C(n1878), .D(n1879), .Y(n1877) );
  XOR2XL U1528 ( .A(\tag_r[4][4] ), .B(proc_addr[9]), .Y(n1878) );
  XOR2XL U1529 ( .A(\tag_r[4][6] ), .B(proc_addr[11]), .Y(n1879) );
  NAND4X1 U1530 ( .A(n1851), .B(n1852), .C(n1853), .D(n1854), .Y(n1850) );
  XOR2XL U1531 ( .A(n1167), .B(proc_addr[26]), .Y(n1853) );
  XOR2XL U1532 ( .A(n1169), .B(proc_addr[24]), .Y(n1852) );
  XOR2XL U1533 ( .A(n1168), .B(proc_addr[25]), .Y(n1851) );
  NAND4X1 U1534 ( .A(n1994), .B(n1995), .C(n1996), .D(n1997), .Y(n1985) );
  XOR2XL U1535 ( .A(n1279), .B(proc_addr[14]), .Y(n1996) );
  XOR2XL U1536 ( .A(n1281), .B(proc_addr[12]), .Y(n1995) );
  XOR2XL U1537 ( .A(n1280), .B(proc_addr[13]), .Y(n1994) );
  NAND4X1 U1538 ( .A(n1858), .B(n1859), .C(n1860), .D(n1861), .Y(n1849) );
  XOR2XL U1539 ( .A(n1179), .B(proc_addr[14]), .Y(n1860) );
  XOR2XL U1540 ( .A(n1181), .B(proc_addr[12]), .Y(n1859) );
  XOR2XL U1541 ( .A(n1180), .B(proc_addr[13]), .Y(n1858) );
  NAND4X1 U1542 ( .A(n1973), .B(n1974), .C(n1975), .D(n1976), .Y(n1946) );
  XOR2XL U1543 ( .A(n1097), .B(proc_addr[21]), .Y(n1975) );
  XOR2XL U1544 ( .A(n1108), .B(proc_addr[10]), .Y(n1974) );
  XOR2XL U1545 ( .A(n1103), .B(proc_addr[15]), .Y(n1973) );
  NAND4X1 U1546 ( .A(n1874), .B(n1875), .C(n1876), .D(n1877), .Y(n1847) );
  XOR2XL U1547 ( .A(n1178), .B(proc_addr[15]), .Y(n1876) );
  XOR2XL U1548 ( .A(n1183), .B(proc_addr[10]), .Y(n1875) );
  XOR2XL U1549 ( .A(n1177), .B(proc_addr[16]), .Y(n1874) );
  NAND4X1 U1550 ( .A(n1866), .B(n1867), .C(n1868), .D(n1869), .Y(n1848) );
  XOR2XL U1551 ( .A(n1165), .B(proc_addr[28]), .Y(n1868) );
  XOR2XL U1552 ( .A(n1166), .B(proc_addr[27]), .Y(n1867) );
  XOR2XL U1553 ( .A(n1164), .B(proc_addr[29]), .Y(n1866) );
  OAI22XL U1554 ( .A0(n4039), .A1(n736), .B0(n1611), .B1(n4032), .Y(n3424) );
  OAI22XL U1555 ( .A0(n4054), .A1(n608), .B0(n1611), .B1(n4045), .Y(n3296) );
  OAI22XL U1556 ( .A0(n4061), .A1(n480), .B0(n1611), .B1(n4064), .Y(n3168) );
  OAI22XL U1557 ( .A0(n4094), .A1(n224), .B0(n1611), .B1(n4088), .Y(n2912) );
  OAI22XL U1558 ( .A0(n4109), .A1(n96), .B0(n1611), .B1(n4102), .Y(n2784) );
  OAI22XL U1559 ( .A0(n4184), .A1(n992), .B0(n1611), .B1(n4178), .Y(n3680) );
  OAI22XL U1560 ( .A0(n4037), .A1(n735), .B0(n1610), .B1(n4035), .Y(n3423) );
  OAI22XL U1561 ( .A0(n4054), .A1(n607), .B0(n1610), .B1(n4044), .Y(n3295) );
  OAI22XL U1562 ( .A0(n4061), .A1(n479), .B0(n1610), .B1(n4064), .Y(n3167) );
  OAI22XL U1563 ( .A0(n4094), .A1(n223), .B0(n1610), .B1(n4088), .Y(n2911) );
  OAI22XL U1564 ( .A0(n4109), .A1(n95), .B0(n1610), .B1(n4102), .Y(n2783) );
  OAI22XL U1565 ( .A0(n4184), .A1(n991), .B0(n1610), .B1(n4177), .Y(n3679) );
  OAI22XL U1566 ( .A0(n4042), .A1(n734), .B0(n1609), .B1(n4032), .Y(n3422) );
  OAI22XL U1567 ( .A0(n4054), .A1(n606), .B0(n1609), .B1(n4047), .Y(n3294) );
  OAI22XL U1568 ( .A0(n4061), .A1(n478), .B0(n1609), .B1(n4064), .Y(n3166) );
  OAI22XL U1569 ( .A0(n4094), .A1(n222), .B0(n1609), .B1(n4088), .Y(n2910) );
  OAI22XL U1570 ( .A0(n4109), .A1(n94), .B0(n1609), .B1(n4102), .Y(n2782) );
  OAI22XL U1571 ( .A0(n1526), .A1(n990), .B0(n1609), .B1(n4183), .Y(n3678) );
  OAI22XL U1572 ( .A0(n4042), .A1(n733), .B0(n1608), .B1(n4033), .Y(n3421) );
  OAI22XL U1573 ( .A0(n4054), .A1(n605), .B0(n1608), .B1(n4044), .Y(n3293) );
  OAI22XL U1574 ( .A0(n4061), .A1(n477), .B0(n1608), .B1(n4064), .Y(n3165) );
  OAI22XL U1575 ( .A0(n4094), .A1(n221), .B0(n1608), .B1(n4088), .Y(n2909) );
  OAI22XL U1576 ( .A0(n4109), .A1(n93), .B0(n1608), .B1(n4102), .Y(n2781) );
  OAI22XL U1577 ( .A0(n1526), .A1(n989), .B0(n1608), .B1(n4178), .Y(n3677) );
  OAI22XL U1578 ( .A0(n4040), .A1(n732), .B0(n1607), .B1(n4029), .Y(n3420) );
  OAI22XL U1579 ( .A0(n4054), .A1(n604), .B0(n1607), .B1(n4043), .Y(n3292) );
  OAI22XL U1580 ( .A0(n4062), .A1(n476), .B0(n1607), .B1(n4064), .Y(n3164) );
  OAI22XL U1581 ( .A0(n4094), .A1(n220), .B0(n1607), .B1(n4088), .Y(n2908) );
  OAI22XL U1582 ( .A0(n4109), .A1(n92), .B0(n1607), .B1(n4102), .Y(n2780) );
  OAI22XL U1583 ( .A0(n1526), .A1(n988), .B0(n1607), .B1(n4177), .Y(n3676) );
  OAI22XL U1584 ( .A0(n4042), .A1(n731), .B0(n1606), .B1(n4033), .Y(n3419) );
  OAI22XL U1585 ( .A0(n4054), .A1(n603), .B0(n1606), .B1(n4047), .Y(n3291) );
  OAI22XL U1586 ( .A0(n4062), .A1(n475), .B0(n1606), .B1(n4064), .Y(n3163) );
  OAI22XL U1587 ( .A0(n4094), .A1(n219), .B0(n1606), .B1(n4088), .Y(n2907) );
  OAI22XL U1588 ( .A0(n4109), .A1(n91), .B0(n1606), .B1(n4102), .Y(n2779) );
  OAI22XL U1589 ( .A0(n1526), .A1(n987), .B0(n1606), .B1(n4183), .Y(n3675) );
  OAI22XL U1590 ( .A0(n4041), .A1(n730), .B0(n1605), .B1(n4035), .Y(n3418) );
  OAI22XL U1591 ( .A0(n4054), .A1(n602), .B0(n1605), .B1(n4044), .Y(n3290) );
  OAI22XL U1592 ( .A0(n4062), .A1(n474), .B0(n1605), .B1(n4064), .Y(n3162) );
  OAI22XL U1593 ( .A0(n4094), .A1(n218), .B0(n1605), .B1(n4088), .Y(n2906) );
  OAI22XL U1594 ( .A0(n4109), .A1(n90), .B0(n1605), .B1(n4102), .Y(n2778) );
  OAI22XL U1595 ( .A0(n4189), .A1(n986), .B0(n1605), .B1(n4181), .Y(n3674) );
  OAI22XL U1596 ( .A0(n4037), .A1(n729), .B0(n1604), .B1(n4032), .Y(n3417) );
  OAI22XL U1597 ( .A0(n4054), .A1(n601), .B0(n1604), .B1(n4047), .Y(n3289) );
  OAI22XL U1598 ( .A0(n4062), .A1(n473), .B0(n1604), .B1(n4067), .Y(n3161) );
  OAI22XL U1599 ( .A0(n4094), .A1(n217), .B0(n1604), .B1(n4088), .Y(n2905) );
  OAI22XL U1600 ( .A0(n4109), .A1(n89), .B0(n1604), .B1(n4102), .Y(n2777) );
  OAI22XL U1601 ( .A0(n4189), .A1(n985), .B0(n1604), .B1(n4181), .Y(n3673) );
  OAI22XL U1602 ( .A0(n4041), .A1(n728), .B0(n1603), .B1(n4033), .Y(n3416) );
  OAI22XL U1603 ( .A0(n4054), .A1(n600), .B0(n1603), .B1(n4044), .Y(n3288) );
  OAI22XL U1604 ( .A0(n4062), .A1(n472), .B0(n1603), .B1(n4068), .Y(n3160) );
  OAI22XL U1605 ( .A0(n4094), .A1(n216), .B0(n1603), .B1(n4088), .Y(n2904) );
  OAI22XL U1606 ( .A0(n4109), .A1(n88), .B0(n1603), .B1(n4102), .Y(n2776) );
  OAI22XL U1607 ( .A0(n4189), .A1(n984), .B0(n1603), .B1(n4181), .Y(n3672) );
  OAI22XL U1608 ( .A0(n4041), .A1(n714), .B0(n1589), .B1(n4034), .Y(n3402) );
  OAI22XL U1609 ( .A0(n4055), .A1(n586), .B0(n1589), .B1(n4048), .Y(n3274) );
  OAI22XL U1610 ( .A0(n4078), .A1(n330), .B0(n1589), .B1(n4073), .Y(n3018) );
  OAI22XL U1611 ( .A0(n4095), .A1(n202), .B0(n1589), .B1(n4089), .Y(n2890) );
  OAI22XL U1612 ( .A0(n4110), .A1(n74), .B0(n1589), .B1(n4103), .Y(n2762) );
  OAI22XL U1613 ( .A0(n4190), .A1(n970), .B0(n1589), .B1(n4182), .Y(n3658) );
  OAI22XL U1614 ( .A0(n4041), .A1(n713), .B0(n1588), .B1(n4034), .Y(n3401) );
  OAI22XL U1615 ( .A0(n4055), .A1(n585), .B0(n1588), .B1(n4048), .Y(n3273) );
  OAI22XL U1616 ( .A0(n4078), .A1(n329), .B0(n1588), .B1(n4073), .Y(n3017) );
  OAI22XL U1617 ( .A0(n4095), .A1(n201), .B0(n1588), .B1(n4089), .Y(n2889) );
  OAI22XL U1618 ( .A0(n4110), .A1(n73), .B0(n1588), .B1(n4103), .Y(n2761) );
  OAI22XL U1619 ( .A0(n4190), .A1(n969), .B0(n1588), .B1(n4182), .Y(n3657) );
  OAI22XL U1620 ( .A0(n4042), .A1(n712), .B0(n1587), .B1(n4034), .Y(n3400) );
  OAI22XL U1621 ( .A0(n4056), .A1(n584), .B0(n1587), .B1(n4046), .Y(n3272) );
  OAI22XL U1622 ( .A0(n4080), .A1(n328), .B0(n1587), .B1(n4072), .Y(n3016) );
  OAI22XL U1623 ( .A0(n4096), .A1(n200), .B0(n1587), .B1(n4083), .Y(n2888) );
  OAI22XL U1624 ( .A0(n4104), .A1(n72), .B0(n1587), .B1(n4097), .Y(n2760) );
  OAI22XL U1625 ( .A0(n4190), .A1(n968), .B0(n1587), .B1(n4182), .Y(n3656) );
  OAI22XL U1626 ( .A0(n4042), .A1(n711), .B0(n1586), .B1(n4034), .Y(n3399) );
  OAI22XL U1627 ( .A0(n4056), .A1(n583), .B0(n1586), .B1(n4048), .Y(n3271) );
  OAI22XL U1628 ( .A0(n4078), .A1(n327), .B0(n1586), .B1(n4073), .Y(n3015) );
  OAI22XL U1629 ( .A0(n4096), .A1(n199), .B0(n1586), .B1(n4089), .Y(n2887) );
  OAI22XL U1630 ( .A0(n4104), .A1(n71), .B0(n1586), .B1(n4103), .Y(n2759) );
  OAI22XL U1631 ( .A0(n4190), .A1(n967), .B0(n1586), .B1(n4182), .Y(n3655) );
  OAI22XL U1632 ( .A0(n1702), .A1(n710), .B0(n1585), .B1(n3), .Y(n3398) );
  OAI22XL U1633 ( .A0(n4056), .A1(n582), .B0(n1585), .B1(n4), .Y(n3270) );
  OAI22XL U1634 ( .A0(n4078), .A1(n326), .B0(n1585), .B1(n4073), .Y(n3014) );
  OAI22XL U1635 ( .A0(n4096), .A1(n198), .B0(n1585), .B1(n4084), .Y(n2886) );
  OAI22XL U1636 ( .A0(n4104), .A1(n70), .B0(n1585), .B1(n4098), .Y(n2758) );
  OAI22XL U1637 ( .A0(n4190), .A1(n966), .B0(n1585), .B1(n4182), .Y(n3654) );
  OAI22XL U1638 ( .A0(n1702), .A1(n709), .B0(n1584), .B1(n3), .Y(n3397) );
  OAI22XL U1639 ( .A0(n4056), .A1(n581), .B0(n1584), .B1(n4), .Y(n3269) );
  OAI22XL U1640 ( .A0(n4078), .A1(n325), .B0(n1584), .B1(n4073), .Y(n3013) );
  OAI22XL U1641 ( .A0(n4096), .A1(n197), .B0(n1584), .B1(n4088), .Y(n2885) );
  OAI22XL U1642 ( .A0(n1578), .A1(n69), .B0(n1584), .B1(n5), .Y(n2757) );
  OAI22XL U1643 ( .A0(n4190), .A1(n965), .B0(n1584), .B1(n4182), .Y(n3653) );
  OAI22XL U1644 ( .A0(n1702), .A1(n708), .B0(n1583), .B1(n3), .Y(n3396) );
  OAI22XL U1645 ( .A0(n4053), .A1(n580), .B0(n1583), .B1(n4), .Y(n3268) );
  OAI22XL U1646 ( .A0(n4080), .A1(n324), .B0(n1583), .B1(n4072), .Y(n3012) );
  OAI22XL U1647 ( .A0(n4096), .A1(n196), .B0(n1583), .B1(n4087), .Y(n2884) );
  OAI22XL U1648 ( .A0(n1578), .A1(n68), .B0(n1583), .B1(n4103), .Y(n2756) );
  OAI22XL U1649 ( .A0(n4190), .A1(n964), .B0(n1583), .B1(n4182), .Y(n3652) );
  OAI22XL U1650 ( .A0(n4042), .A1(n707), .B0(n1582), .B1(n3), .Y(n3395) );
  OAI22XL U1651 ( .A0(n4055), .A1(n579), .B0(n1582), .B1(n4), .Y(n3267) );
  OAI22XL U1652 ( .A0(n1694), .A1(n323), .B0(n1582), .B1(n4073), .Y(n3011) );
  OAI22XL U1653 ( .A0(n4096), .A1(n195), .B0(n1582), .B1(n4085), .Y(n2883) );
  OAI22XL U1654 ( .A0(n1578), .A1(n67), .B0(n1582), .B1(n5), .Y(n2755) );
  OAI22XL U1655 ( .A0(n4190), .A1(n963), .B0(n1582), .B1(n4182), .Y(n3651) );
  OAI22XL U1656 ( .A0(n4042), .A1(n706), .B0(n1581), .B1(n4030), .Y(n3394) );
  OAI22XL U1657 ( .A0(n4056), .A1(n578), .B0(n1581), .B1(n4045), .Y(n3266) );
  OAI22XL U1658 ( .A0(n4081), .A1(n322), .B0(n1581), .B1(n4072), .Y(n3010) );
  OAI22XL U1659 ( .A0(n4096), .A1(n194), .B0(n1581), .B1(n4087), .Y(n2882) );
  OAI22XL U1660 ( .A0(n4104), .A1(n66), .B0(n1581), .B1(n4100), .Y(n2754) );
  OAI22XL U1661 ( .A0(n4187), .A1(n962), .B0(n1581), .B1(n4183), .Y(n3650) );
  OAI22XL U1662 ( .A0(n4042), .A1(n705), .B0(n1579), .B1(n4031), .Y(n3393) );
  OAI22XL U1663 ( .A0(n4056), .A1(n577), .B0(n1579), .B1(n4046), .Y(n3265) );
  OAI22XL U1664 ( .A0(n1694), .A1(n321), .B0(n1579), .B1(n4074), .Y(n3009) );
  OAI22XL U1665 ( .A0(n4096), .A1(n193), .B0(n1579), .B1(n4086), .Y(n2881) );
  OAI22XL U1666 ( .A0(n1578), .A1(n65), .B0(n1579), .B1(n4102), .Y(n2753) );
  OAI22XL U1667 ( .A0(n4188), .A1(n961), .B0(n1579), .B1(n4183), .Y(n3649) );
  OAI22XL U1668 ( .A0(n4037), .A1(n813), .B0(n1688), .B1(n4029), .Y(n3501) );
  OAI22XL U1669 ( .A0(n4053), .A1(n685), .B0(n1688), .B1(n4043), .Y(n3373) );
  OAI22XL U1670 ( .A0(n4079), .A1(n429), .B0(n1688), .B1(n4076), .Y(n3117) );
  OAI22XL U1671 ( .A0(n4091), .A1(n301), .B0(n1688), .B1(n4084), .Y(n2989) );
  OAI22XL U1672 ( .A0(n4106), .A1(n173), .B0(n1688), .B1(n4098), .Y(n2861) );
  OAI22XL U1673 ( .A0(n4190), .A1(n1069), .B0(n1688), .B1(n4177), .Y(n3757) );
  OAI22XL U1674 ( .A0(n4040), .A1(n812), .B0(n1687), .B1(n4029), .Y(n3500) );
  OAI22XL U1675 ( .A0(n4055), .A1(n684), .B0(n1687), .B1(n4043), .Y(n3372) );
  OAI22XL U1676 ( .A0(n4079), .A1(n428), .B0(n1687), .B1(n4076), .Y(n3116) );
  OAI22XL U1677 ( .A0(n4092), .A1(n300), .B0(n1687), .B1(n4084), .Y(n2988) );
  OAI22XL U1678 ( .A0(n4110), .A1(n172), .B0(n1687), .B1(n4098), .Y(n2860) );
  OAI22XL U1679 ( .A0(n4189), .A1(n1068), .B0(n1687), .B1(n4177), .Y(n3756) );
  OAI22XL U1680 ( .A0(n4041), .A1(n811), .B0(n1686), .B1(n4029), .Y(n3499) );
  OAI22XL U1681 ( .A0(n4051), .A1(n683), .B0(n1686), .B1(n4043), .Y(n3371) );
  OAI22XL U1682 ( .A0(n4079), .A1(n427), .B0(n1686), .B1(n4076), .Y(n3115) );
  OAI22XL U1683 ( .A0(n4095), .A1(n299), .B0(n1686), .B1(n4084), .Y(n2987) );
  OAI22XL U1684 ( .A0(n4110), .A1(n171), .B0(n1686), .B1(n4098), .Y(n2859) );
  OAI22XL U1685 ( .A0(n4186), .A1(n1067), .B0(n1686), .B1(n4177), .Y(n3755) );
  OAI22XL U1686 ( .A0(n4039), .A1(n810), .B0(n1685), .B1(n4029), .Y(n3498) );
  OAI22XL U1687 ( .A0(n4050), .A1(n682), .B0(n1685), .B1(n4043), .Y(n3370) );
  OAI22XL U1688 ( .A0(n4079), .A1(n426), .B0(n1685), .B1(n4076), .Y(n3114) );
  OAI22XL U1689 ( .A0(n4096), .A1(n298), .B0(n1685), .B1(n4084), .Y(n2986) );
  OAI22XL U1690 ( .A0(n4107), .A1(n170), .B0(n1685), .B1(n4098), .Y(n2858) );
  OAI22XL U1691 ( .A0(n4185), .A1(n1066), .B0(n1685), .B1(n4177), .Y(n3754) );
  OAI22XL U1692 ( .A0(n4038), .A1(n809), .B0(n1684), .B1(n4029), .Y(n3497) );
  OAI22XL U1693 ( .A0(n4050), .A1(n681), .B0(n1684), .B1(n4043), .Y(n3369) );
  OAI22XL U1694 ( .A0(n4079), .A1(n425), .B0(n1684), .B1(n4076), .Y(n3113) );
  OAI22XL U1695 ( .A0(n4092), .A1(n297), .B0(n1684), .B1(n4084), .Y(n2985) );
  OAI22XL U1696 ( .A0(n4108), .A1(n169), .B0(n1684), .B1(n4098), .Y(n2857) );
  OAI22XL U1697 ( .A0(n4184), .A1(n1065), .B0(n1684), .B1(n4177), .Y(n3753) );
  OAI22XL U1698 ( .A0(n4036), .A1(n808), .B0(n1683), .B1(n4035), .Y(n3496) );
  OAI22XL U1699 ( .A0(n4050), .A1(n680), .B0(n1683), .B1(n4044), .Y(n3368) );
  OAI22XL U1700 ( .A0(n4079), .A1(n424), .B0(n1683), .B1(n4076), .Y(n3112) );
  OAI22XL U1701 ( .A0(n4091), .A1(n296), .B0(n1683), .B1(n4085), .Y(n2984) );
  OAI22XL U1702 ( .A0(n4105), .A1(n168), .B0(n1683), .B1(n4099), .Y(n2856) );
  OAI22XL U1703 ( .A0(n4185), .A1(n1064), .B0(n1683), .B1(n4177), .Y(n3752) );
  OAI22XL U1704 ( .A0(n4036), .A1(n807), .B0(n1682), .B1(n4035), .Y(n3495) );
  OAI22XL U1705 ( .A0(n4050), .A1(n679), .B0(n1682), .B1(n4044), .Y(n3367) );
  OAI22XL U1706 ( .A0(n4079), .A1(n423), .B0(n1682), .B1(n4076), .Y(n3111) );
  OAI22XL U1707 ( .A0(n4091), .A1(n295), .B0(n1682), .B1(n4085), .Y(n2983) );
  OAI22XL U1708 ( .A0(n4105), .A1(n167), .B0(n1682), .B1(n4099), .Y(n2855) );
  OAI22XL U1709 ( .A0(n4184), .A1(n1063), .B0(n1682), .B1(n4177), .Y(n3751) );
  OAI22XL U1710 ( .A0(n4036), .A1(n806), .B0(n1681), .B1(n4035), .Y(n3494) );
  OAI22XL U1711 ( .A0(n4050), .A1(n678), .B0(n1681), .B1(n4044), .Y(n3366) );
  OAI22XL U1712 ( .A0(n4079), .A1(n422), .B0(n1681), .B1(n4076), .Y(n3110) );
  OAI22XL U1713 ( .A0(n4091), .A1(n294), .B0(n1681), .B1(n4085), .Y(n2982) );
  OAI22XL U1714 ( .A0(n4105), .A1(n166), .B0(n1681), .B1(n4099), .Y(n2854) );
  OAI22XL U1715 ( .A0(n4190), .A1(n1062), .B0(n1681), .B1(n4177), .Y(n3750) );
  OAI22XL U1716 ( .A0(n4036), .A1(n805), .B0(n1680), .B1(n4035), .Y(n3493) );
  OAI22XL U1717 ( .A0(n4050), .A1(n677), .B0(n1680), .B1(n4044), .Y(n3365) );
  OAI22XL U1718 ( .A0(n4079), .A1(n421), .B0(n1680), .B1(n4076), .Y(n3109) );
  OAI22XL U1719 ( .A0(n4091), .A1(n293), .B0(n1680), .B1(n4085), .Y(n2981) );
  OAI22XL U1720 ( .A0(n4105), .A1(n165), .B0(n1680), .B1(n4099), .Y(n2853) );
  OAI22XL U1721 ( .A0(n4189), .A1(n1061), .B0(n1680), .B1(n4177), .Y(n3749) );
  OAI22XL U1722 ( .A0(n4036), .A1(n804), .B0(n1679), .B1(n4035), .Y(n3492) );
  OAI22XL U1723 ( .A0(n4050), .A1(n676), .B0(n1679), .B1(n4044), .Y(n3364) );
  OAI22XL U1724 ( .A0(n4079), .A1(n420), .B0(n1679), .B1(n4076), .Y(n3108) );
  OAI22XL U1725 ( .A0(n4091), .A1(n292), .B0(n1679), .B1(n4085), .Y(n2980) );
  OAI22XL U1726 ( .A0(n4105), .A1(n164), .B0(n1679), .B1(n4099), .Y(n2852) );
  OAI22XL U1727 ( .A0(n4190), .A1(n1060), .B0(n1679), .B1(n4177), .Y(n3748) );
  OAI22XL U1728 ( .A0(n4036), .A1(n803), .B0(n1678), .B1(n4035), .Y(n3491) );
  OAI22XL U1729 ( .A0(n4050), .A1(n675), .B0(n1678), .B1(n4044), .Y(n3363) );
  OAI22XL U1730 ( .A0(n4079), .A1(n419), .B0(n1678), .B1(n4076), .Y(n3107) );
  OAI22XL U1731 ( .A0(n4091), .A1(n291), .B0(n1678), .B1(n4085), .Y(n2979) );
  OAI22XL U1732 ( .A0(n4105), .A1(n163), .B0(n1678), .B1(n4099), .Y(n2851) );
  OAI22XL U1733 ( .A0(n4185), .A1(n1059), .B0(n1678), .B1(n4177), .Y(n3747) );
  OAI22XL U1734 ( .A0(n4036), .A1(n802), .B0(n1677), .B1(n4035), .Y(n3490) );
  OAI22XL U1735 ( .A0(n4050), .A1(n674), .B0(n1677), .B1(n4044), .Y(n3362) );
  OAI22XL U1736 ( .A0(n4080), .A1(n418), .B0(n1677), .B1(n4076), .Y(n3106) );
  OAI22XL U1737 ( .A0(n4091), .A1(n290), .B0(n1677), .B1(n4085), .Y(n2978) );
  OAI22XL U1738 ( .A0(n4105), .A1(n162), .B0(n1677), .B1(n4099), .Y(n2850) );
  OAI22XL U1739 ( .A0(n4185), .A1(n1058), .B0(n1677), .B1(n4178), .Y(n3746) );
  OAI22XL U1740 ( .A0(n4036), .A1(n801), .B0(n1676), .B1(n4035), .Y(n3489) );
  OAI22XL U1741 ( .A0(n4050), .A1(n673), .B0(n1676), .B1(n4044), .Y(n3361) );
  OAI22XL U1742 ( .A0(n4080), .A1(n417), .B0(n1676), .B1(n4076), .Y(n3105) );
  OAI22XL U1743 ( .A0(n4091), .A1(n289), .B0(n1676), .B1(n4085), .Y(n2977) );
  OAI22XL U1744 ( .A0(n4105), .A1(n161), .B0(n1676), .B1(n4099), .Y(n2849) );
  OAI22XL U1745 ( .A0(n4185), .A1(n1057), .B0(n1676), .B1(n4178), .Y(n3745) );
  OAI22XL U1746 ( .A0(n4036), .A1(n800), .B0(n1675), .B1(n4035), .Y(n3488) );
  OAI22XL U1747 ( .A0(n4050), .A1(n672), .B0(n1675), .B1(n4044), .Y(n3360) );
  OAI22XL U1748 ( .A0(n4080), .A1(n416), .B0(n1675), .B1(n4076), .Y(n3104) );
  OAI22XL U1749 ( .A0(n4091), .A1(n288), .B0(n1675), .B1(n4085), .Y(n2976) );
  OAI22XL U1750 ( .A0(n4105), .A1(n160), .B0(n1675), .B1(n4099), .Y(n2848) );
  OAI22XL U1751 ( .A0(n4185), .A1(n1056), .B0(n1675), .B1(n4178), .Y(n3744) );
  OAI22XL U1752 ( .A0(n4036), .A1(n799), .B0(n1674), .B1(n4034), .Y(n3487) );
  OAI22XL U1753 ( .A0(n4050), .A1(n671), .B0(n1674), .B1(n4044), .Y(n3359) );
  OAI22XL U1754 ( .A0(n4080), .A1(n415), .B0(n1674), .B1(n4076), .Y(n3103) );
  OAI22XL U1755 ( .A0(n4091), .A1(n287), .B0(n1674), .B1(n4085), .Y(n2975) );
  OAI22XL U1756 ( .A0(n4105), .A1(n159), .B0(n1674), .B1(n4099), .Y(n2847) );
  OAI22XL U1757 ( .A0(n4185), .A1(n1055), .B0(n1674), .B1(n4178), .Y(n3743) );
  OAI22XL U1758 ( .A0(n4036), .A1(n798), .B0(n1673), .B1(n4031), .Y(n3486) );
  OAI22XL U1759 ( .A0(n4050), .A1(n670), .B0(n1673), .B1(n4044), .Y(n3358) );
  OAI22XL U1760 ( .A0(n4080), .A1(n414), .B0(n1673), .B1(n4075), .Y(n3102) );
  OAI22XL U1761 ( .A0(n4091), .A1(n286), .B0(n1673), .B1(n4085), .Y(n2974) );
  OAI22XL U1762 ( .A0(n4105), .A1(n158), .B0(n1673), .B1(n4099), .Y(n2846) );
  OAI22XL U1763 ( .A0(n4185), .A1(n1054), .B0(n1673), .B1(n4178), .Y(n3742) );
  OAI22XL U1764 ( .A0(n4041), .A1(n743), .B0(n1618), .B1(n4030), .Y(n3431) );
  OAI22XL U1765 ( .A0(n4053), .A1(n615), .B0(n1618), .B1(n4048), .Y(n3303) );
  OAI22XL U1766 ( .A0(n4061), .A1(n487), .B0(n1618), .B1(n4065), .Y(n3175) );
  OAI22XL U1767 ( .A0(n4096), .A1(n231), .B0(n1618), .B1(n4087), .Y(n2919) );
  OAI22XL U1768 ( .A0(n4107), .A1(n103), .B0(n1618), .B1(n4102), .Y(n2791) );
  OAI22XL U1769 ( .A0(n4187), .A1(n999), .B0(n1618), .B1(n4178), .Y(n3687) );
  OAI22XL U1770 ( .A0(n4037), .A1(n742), .B0(n1617), .B1(n4032), .Y(n3430) );
  OAI22XL U1771 ( .A0(n4053), .A1(n614), .B0(n1617), .B1(n4045), .Y(n3302) );
  OAI22XL U1772 ( .A0(n4061), .A1(n486), .B0(n1617), .B1(n4065), .Y(n3174) );
  OAI22XL U1773 ( .A0(n4096), .A1(n230), .B0(n1617), .B1(n4087), .Y(n2918) );
  OAI22XL U1774 ( .A0(n4108), .A1(n102), .B0(n1617), .B1(n4103), .Y(n2790) );
  OAI22XL U1775 ( .A0(n1526), .A1(n998), .B0(n1617), .B1(n4178), .Y(n3686) );
  OAI22XL U1776 ( .A0(n4041), .A1(n741), .B0(n1616), .B1(n4033), .Y(n3429) );
  OAI22XL U1777 ( .A0(n4053), .A1(n613), .B0(n1616), .B1(n4047), .Y(n3301) );
  OAI22XL U1778 ( .A0(n4061), .A1(n485), .B0(n1616), .B1(n4065), .Y(n3173) );
  OAI22XL U1779 ( .A0(n4096), .A1(n229), .B0(n1616), .B1(n4087), .Y(n2917) );
  OAI22XL U1780 ( .A0(n4107), .A1(n101), .B0(n1616), .B1(n4102), .Y(n2789) );
  OAI22XL U1781 ( .A0(n4184), .A1(n997), .B0(n1616), .B1(n4177), .Y(n3685) );
  OAI22XL U1782 ( .A0(n4041), .A1(n740), .B0(n1615), .B1(n4034), .Y(n3428) );
  OAI22XL U1783 ( .A0(n4053), .A1(n612), .B0(n1615), .B1(n4046), .Y(n3300) );
  OAI22XL U1784 ( .A0(n4061), .A1(n484), .B0(n1615), .B1(n4065), .Y(n3172) );
  OAI22XL U1785 ( .A0(n4096), .A1(n228), .B0(n1615), .B1(n4087), .Y(n2916) );
  OAI22XL U1786 ( .A0(n4109), .A1(n100), .B0(n1615), .B1(n4103), .Y(n2788) );
  OAI22XL U1787 ( .A0(n4184), .A1(n996), .B0(n1615), .B1(n4183), .Y(n3684) );
  OAI22XL U1788 ( .A0(n4037), .A1(n739), .B0(n1614), .B1(n4031), .Y(n3427) );
  OAI22XL U1789 ( .A0(n4053), .A1(n611), .B0(n1614), .B1(n4043), .Y(n3299) );
  OAI22XL U1790 ( .A0(n4061), .A1(n483), .B0(n1614), .B1(n4065), .Y(n3171) );
  OAI22XL U1791 ( .A0(n4092), .A1(n227), .B0(n1614), .B1(n4087), .Y(n2915) );
  OAI22XL U1792 ( .A0(n4105), .A1(n99), .B0(n1614), .B1(n4102), .Y(n2787) );
  OAI22XL U1793 ( .A0(n4184), .A1(n995), .B0(n1614), .B1(n4178), .Y(n3683) );
  OAI22XL U1794 ( .A0(n4040), .A1(n738), .B0(n1613), .B1(n4029), .Y(n3426) );
  OAI22XL U1795 ( .A0(n4053), .A1(n610), .B0(n1613), .B1(n4044), .Y(n3298) );
  OAI22XL U1796 ( .A0(n4061), .A1(n482), .B0(n1613), .B1(n4067), .Y(n3170) );
  OAI22XL U1797 ( .A0(n4095), .A1(n226), .B0(n1613), .B1(n4087), .Y(n2914) );
  OAI22XL U1798 ( .A0(n4104), .A1(n98), .B0(n1613), .B1(n4103), .Y(n2786) );
  OAI22XL U1799 ( .A0(n4184), .A1(n994), .B0(n1613), .B1(n4177), .Y(n3682) );
  OAI22XL U1800 ( .A0(n4039), .A1(n737), .B0(n1612), .B1(n4035), .Y(n3425) );
  OAI22XL U1801 ( .A0(n4053), .A1(n609), .B0(n1612), .B1(n4049), .Y(n3297) );
  OAI22XL U1802 ( .A0(n4061), .A1(n481), .B0(n1612), .B1(n4066), .Y(n3169) );
  OAI22XL U1803 ( .A0(n4096), .A1(n225), .B0(n1612), .B1(n4087), .Y(n2913) );
  OAI22XL U1804 ( .A0(n4104), .A1(n97), .B0(n1612), .B1(n4102), .Y(n2785) );
  OAI22XL U1805 ( .A0(n4184), .A1(n993), .B0(n1612), .B1(n4183), .Y(n3681) );
  OAI22XL U1806 ( .A0(n4039), .A1(n832), .B0(n1545), .B1(n4031), .Y(n3520) );
  OAI22XL U1807 ( .A0(n4052), .A1(n704), .B0(n1545), .B1(n4048), .Y(n3392) );
  OAI22XL U1808 ( .A0(n4062), .A1(n576), .B0(n1545), .B1(n4068), .Y(n3264) );
  OAI22XL U1809 ( .A0(n4093), .A1(n320), .B0(n1545), .B1(n4083), .Y(n3008) );
  OAI22XL U1810 ( .A0(n4106), .A1(n192), .B0(n1545), .B1(n4097), .Y(n2880) );
  OAI22XL U1811 ( .A0(n4184), .A1(n1088), .B0(n1545), .B1(n4183), .Y(n3776) );
  OAI22XL U1812 ( .A0(n4036), .A1(n831), .B0(n1544), .B1(n4030), .Y(n3519) );
  OAI22XL U1813 ( .A0(n4056), .A1(n703), .B0(n1544), .B1(n4045), .Y(n3391) );
  OAI22XL U1814 ( .A0(n4059), .A1(n575), .B0(n1544), .B1(n4070), .Y(n3263) );
  OAI22XL U1815 ( .A0(n4090), .A1(n319), .B0(n1544), .B1(n4083), .Y(n3007) );
  OAI22XL U1816 ( .A0(n4106), .A1(n191), .B0(n1544), .B1(n4097), .Y(n2879) );
  OAI22XL U1817 ( .A0(n4184), .A1(n1087), .B0(n1544), .B1(n4183), .Y(n3775) );
  OAI22XL U1818 ( .A0(n4040), .A1(n830), .B0(n1543), .B1(n4034), .Y(n3518) );
  OAI22XL U1819 ( .A0(n4052), .A1(n702), .B0(n1543), .B1(n4046), .Y(n3390) );
  OAI22XL U1820 ( .A0(n4057), .A1(n574), .B0(n1543), .B1(n4070), .Y(n3262) );
  OAI22XL U1821 ( .A0(n4094), .A1(n318), .B0(n1543), .B1(n4083), .Y(n3006) );
  OAI22XL U1822 ( .A0(n4110), .A1(n190), .B0(n1543), .B1(n4097), .Y(n2878) );
  OAI22XL U1823 ( .A0(n4184), .A1(n1086), .B0(n1543), .B1(n4183), .Y(n3774) );
  OAI22XL U1824 ( .A0(n4038), .A1(n829), .B0(n1542), .B1(n4031), .Y(n3517) );
  OAI22XL U1825 ( .A0(n4054), .A1(n701), .B0(n1542), .B1(n4048), .Y(n3389) );
  OAI22XL U1826 ( .A0(n4057), .A1(n573), .B0(n1542), .B1(n4070), .Y(n3261) );
  OAI22XL U1827 ( .A0(n4094), .A1(n317), .B0(n1542), .B1(n4083), .Y(n3005) );
  OAI22XL U1828 ( .A0(n4107), .A1(n189), .B0(n1542), .B1(n4097), .Y(n2877) );
  OAI22XL U1829 ( .A0(n4184), .A1(n1085), .B0(n1542), .B1(n4183), .Y(n3773) );
  OAI22XL U1830 ( .A0(n4039), .A1(n828), .B0(n1541), .B1(n4030), .Y(n3516) );
  OAI22XL U1831 ( .A0(n4056), .A1(n700), .B0(n1541), .B1(n4045), .Y(n3388) );
  OAI22XL U1832 ( .A0(n4062), .A1(n572), .B0(n1541), .B1(n4070), .Y(n3260) );
  OAI22XL U1833 ( .A0(n4091), .A1(n316), .B0(n1541), .B1(n4083), .Y(n3004) );
  OAI22XL U1834 ( .A0(n4108), .A1(n188), .B0(n1541), .B1(n4097), .Y(n2876) );
  OAI22XL U1835 ( .A0(n4185), .A1(n1084), .B0(n1541), .B1(n4183), .Y(n3772) );
  OAI22XL U1836 ( .A0(n4037), .A1(n827), .B0(n1540), .B1(n4029), .Y(n3515) );
  OAI22XL U1837 ( .A0(n4052), .A1(n699), .B0(n1540), .B1(n4043), .Y(n3387) );
  OAI22XL U1838 ( .A0(n4061), .A1(n571), .B0(n1540), .B1(n4070), .Y(n3259) );
  OAI22XL U1839 ( .A0(n4091), .A1(n315), .B0(n1540), .B1(n4083), .Y(n3003) );
  OAI22XL U1840 ( .A0(n4109), .A1(n187), .B0(n1540), .B1(n4097), .Y(n2875) );
  OAI22XL U1841 ( .A0(n4186), .A1(n1083), .B0(n1540), .B1(n4183), .Y(n3771) );
  OAI22XL U1842 ( .A0(n4036), .A1(n727), .B0(n1602), .B1(n4029), .Y(n3415) );
  OAI22XL U1843 ( .A0(n4054), .A1(n599), .B0(n1602), .B1(n4043), .Y(n3287) );
  OAI22XL U1844 ( .A0(n4062), .A1(n471), .B0(n1602), .B1(n4064), .Y(n3159) );
  OAI22XL U1845 ( .A0(n4080), .A1(n343), .B0(n1602), .B1(n4077), .Y(n3031) );
  OAI22XL U1846 ( .A0(n4094), .A1(n215), .B0(n1602), .B1(n4088), .Y(n2903) );
  OAI22XL U1847 ( .A0(n4109), .A1(n87), .B0(n1602), .B1(n4102), .Y(n2775) );
  OAI22XL U1848 ( .A0(n4189), .A1(n983), .B0(n1602), .B1(n4181), .Y(n3671) );
  OAI22XL U1849 ( .A0(n4038), .A1(n726), .B0(n1601), .B1(n4035), .Y(n3414) );
  OAI22XL U1850 ( .A0(n4054), .A1(n598), .B0(n1601), .B1(n4049), .Y(n3286) );
  OAI22XL U1851 ( .A0(n4062), .A1(n470), .B0(n1601), .B1(n4067), .Y(n3158) );
  OAI22XL U1852 ( .A0(n4082), .A1(n342), .B0(n1601), .B1(n4077), .Y(n3030) );
  OAI22XL U1853 ( .A0(n4094), .A1(n214), .B0(n1601), .B1(n4088), .Y(n2902) );
  OAI22XL U1854 ( .A0(n4109), .A1(n86), .B0(n1601), .B1(n4102), .Y(n2774) );
  OAI22XL U1855 ( .A0(n4189), .A1(n982), .B0(n1601), .B1(n4181), .Y(n3670) );
  OAI22XL U1856 ( .A0(n4039), .A1(n725), .B0(n1600), .B1(n3), .Y(n3413) );
  OAI22XL U1857 ( .A0(n4054), .A1(n597), .B0(n1600), .B1(n4), .Y(n3285) );
  OAI22XL U1858 ( .A0(n4062), .A1(n469), .B0(n1600), .B1(n4068), .Y(n3157) );
  OAI22XL U1859 ( .A0(n4082), .A1(n341), .B0(n1600), .B1(n4073), .Y(n3029) );
  OAI22XL U1860 ( .A0(n4094), .A1(n213), .B0(n1600), .B1(n4088), .Y(n2901) );
  OAI22XL U1861 ( .A0(n4109), .A1(n85), .B0(n1600), .B1(n4102), .Y(n2773) );
  OAI22XL U1862 ( .A0(n4189), .A1(n981), .B0(n1600), .B1(n4181), .Y(n3669) );
  OAI22XL U1863 ( .A0(n4041), .A1(n724), .B0(n1599), .B1(n4034), .Y(n3412) );
  OAI22XL U1864 ( .A0(n4055), .A1(n596), .B0(n1599), .B1(n4048), .Y(n3284) );
  OAI22XL U1865 ( .A0(n4062), .A1(n468), .B0(n1599), .B1(n4067), .Y(n3156) );
  OAI22XL U1866 ( .A0(n4082), .A1(n340), .B0(n1599), .B1(n4073), .Y(n3028) );
  OAI22XL U1867 ( .A0(n4095), .A1(n212), .B0(n1599), .B1(n4089), .Y(n2900) );
  OAI22XL U1868 ( .A0(n4110), .A1(n84), .B0(n1599), .B1(n4103), .Y(n2772) );
  OAI22XL U1869 ( .A0(n4189), .A1(n980), .B0(n1599), .B1(n4181), .Y(n3668) );
  OAI22XL U1870 ( .A0(n4041), .A1(n723), .B0(n1598), .B1(n4034), .Y(n3411) );
  OAI22XL U1871 ( .A0(n4055), .A1(n595), .B0(n1598), .B1(n4048), .Y(n3283) );
  OAI22XL U1872 ( .A0(n4062), .A1(n467), .B0(n1598), .B1(n4068), .Y(n3155) );
  OAI22XL U1873 ( .A0(n4082), .A1(n339), .B0(n1598), .B1(n4072), .Y(n3027) );
  OAI22XL U1874 ( .A0(n4095), .A1(n211), .B0(n1598), .B1(n4089), .Y(n2899) );
  OAI22XL U1875 ( .A0(n4110), .A1(n83), .B0(n1598), .B1(n4103), .Y(n2771) );
  OAI22XL U1876 ( .A0(n4189), .A1(n979), .B0(n1598), .B1(n4181), .Y(n3667) );
  OAI22XL U1877 ( .A0(n4041), .A1(n722), .B0(n1597), .B1(n4034), .Y(n3410) );
  OAI22XL U1878 ( .A0(n4055), .A1(n594), .B0(n1597), .B1(n4048), .Y(n3282) );
  OAI22XL U1879 ( .A0(n4062), .A1(n466), .B0(n1597), .B1(n4064), .Y(n3154) );
  OAI22XL U1880 ( .A0(n4082), .A1(n338), .B0(n1597), .B1(n4073), .Y(n3026) );
  OAI22XL U1881 ( .A0(n4095), .A1(n210), .B0(n1597), .B1(n4089), .Y(n2898) );
  OAI22XL U1882 ( .A0(n4110), .A1(n82), .B0(n1597), .B1(n4103), .Y(n2770) );
  OAI22XL U1883 ( .A0(n4189), .A1(n978), .B0(n1597), .B1(n4181), .Y(n3666) );
  OAI22XL U1884 ( .A0(n4041), .A1(n721), .B0(n1596), .B1(n4034), .Y(n3409) );
  OAI22XL U1885 ( .A0(n4055), .A1(n593), .B0(n1596), .B1(n4048), .Y(n3281) );
  OAI22XL U1886 ( .A0(n4062), .A1(n465), .B0(n1596), .B1(n4065), .Y(n3153) );
  OAI22XL U1887 ( .A0(n4082), .A1(n337), .B0(n1596), .B1(n4077), .Y(n3025) );
  OAI22XL U1888 ( .A0(n4095), .A1(n209), .B0(n1596), .B1(n4089), .Y(n2897) );
  OAI22XL U1889 ( .A0(n4110), .A1(n81), .B0(n1596), .B1(n4103), .Y(n2769) );
  OAI22XL U1890 ( .A0(n4189), .A1(n977), .B0(n1596), .B1(n4181), .Y(n3665) );
  OAI22XL U1891 ( .A0(n4041), .A1(n720), .B0(n1595), .B1(n4034), .Y(n3408) );
  OAI22XL U1892 ( .A0(n4055), .A1(n592), .B0(n1595), .B1(n4048), .Y(n3280) );
  OAI22XL U1893 ( .A0(n4060), .A1(n464), .B0(n1595), .B1(n4066), .Y(n3152) );
  OAI22XL U1894 ( .A0(n4082), .A1(n336), .B0(n1595), .B1(n4073), .Y(n3024) );
  OAI22XL U1895 ( .A0(n4095), .A1(n208), .B0(n1595), .B1(n4089), .Y(n2896) );
  OAI22XL U1896 ( .A0(n4110), .A1(n80), .B0(n1595), .B1(n4103), .Y(n2768) );
  OAI22XL U1897 ( .A0(n4189), .A1(n976), .B0(n1595), .B1(n4181), .Y(n3664) );
  OAI22XL U1898 ( .A0(n4041), .A1(n719), .B0(n1594), .B1(n4034), .Y(n3407) );
  OAI22XL U1899 ( .A0(n4055), .A1(n591), .B0(n1594), .B1(n4048), .Y(n3279) );
  OAI22XL U1900 ( .A0(n4062), .A1(n463), .B0(n1594), .B1(n8), .Y(n3151) );
  OAI22XL U1901 ( .A0(n4082), .A1(n335), .B0(n1594), .B1(n4073), .Y(n3023) );
  OAI22XL U1902 ( .A0(n4095), .A1(n207), .B0(n1594), .B1(n4089), .Y(n2895) );
  OAI22XL U1903 ( .A0(n4110), .A1(n79), .B0(n1594), .B1(n4103), .Y(n2767) );
  OAI22XL U1904 ( .A0(n4189), .A1(n975), .B0(n1594), .B1(n4181), .Y(n3663) );
  OAI22XL U1905 ( .A0(n4041), .A1(n718), .B0(n1593), .B1(n4034), .Y(n3406) );
  OAI22XL U1906 ( .A0(n4055), .A1(n590), .B0(n1593), .B1(n4048), .Y(n3278) );
  OAI22XL U1907 ( .A0(n4058), .A1(n462), .B0(n1593), .B1(n4065), .Y(n3150) );
  OAI22XL U1908 ( .A0(n4082), .A1(n334), .B0(n1593), .B1(n4073), .Y(n3022) );
  OAI22XL U1909 ( .A0(n4095), .A1(n206), .B0(n1593), .B1(n4089), .Y(n2894) );
  OAI22XL U1910 ( .A0(n4110), .A1(n78), .B0(n1593), .B1(n4103), .Y(n2766) );
  OAI22XL U1911 ( .A0(n4190), .A1(n974), .B0(n1593), .B1(n4182), .Y(n3662) );
  OAI22XL U1912 ( .A0(n4041), .A1(n717), .B0(n1592), .B1(n4034), .Y(n3405) );
  OAI22XL U1913 ( .A0(n4055), .A1(n589), .B0(n1592), .B1(n4048), .Y(n3277) );
  OAI22XL U1914 ( .A0(n4059), .A1(n461), .B0(n1592), .B1(n4066), .Y(n3149) );
  OAI22XL U1915 ( .A0(n4082), .A1(n333), .B0(n1592), .B1(n4073), .Y(n3021) );
  OAI22XL U1916 ( .A0(n4095), .A1(n205), .B0(n1592), .B1(n4089), .Y(n2893) );
  OAI22XL U1917 ( .A0(n4110), .A1(n77), .B0(n1592), .B1(n4103), .Y(n2765) );
  OAI22XL U1918 ( .A0(n4190), .A1(n973), .B0(n1592), .B1(n4182), .Y(n3661) );
  OAI22XL U1919 ( .A0(n4041), .A1(n716), .B0(n1591), .B1(n4034), .Y(n3404) );
  OAI22XL U1920 ( .A0(n4055), .A1(n588), .B0(n1591), .B1(n4048), .Y(n3276) );
  OAI22XL U1921 ( .A0(n4061), .A1(n460), .B0(n1591), .B1(n4065), .Y(n3148) );
  OAI22XL U1922 ( .A0(n4082), .A1(n332), .B0(n1591), .B1(n4073), .Y(n3020) );
  OAI22XL U1923 ( .A0(n4095), .A1(n204), .B0(n1591), .B1(n4089), .Y(n2892) );
  OAI22XL U1924 ( .A0(n4110), .A1(n76), .B0(n1591), .B1(n4103), .Y(n2764) );
  OAI22XL U1925 ( .A0(n4190), .A1(n972), .B0(n1591), .B1(n4182), .Y(n3660) );
  OAI22XL U1926 ( .A0(n4041), .A1(n715), .B0(n1590), .B1(n4034), .Y(n3403) );
  OAI22XL U1927 ( .A0(n4055), .A1(n587), .B0(n1590), .B1(n4048), .Y(n3275) );
  OAI22XL U1928 ( .A0(n4060), .A1(n459), .B0(n1590), .B1(n4066), .Y(n3147) );
  OAI22XL U1929 ( .A0(n4082), .A1(n331), .B0(n1590), .B1(n4073), .Y(n3019) );
  OAI22XL U1930 ( .A0(n4095), .A1(n203), .B0(n1590), .B1(n4089), .Y(n2891) );
  OAI22XL U1931 ( .A0(n4110), .A1(n75), .B0(n1590), .B1(n4103), .Y(n2763) );
  OAI22XL U1932 ( .A0(n4190), .A1(n971), .B0(n1590), .B1(n4182), .Y(n3659) );
  OAI22XL U1933 ( .A0(n4036), .A1(n814), .B0(n1689), .B1(n4029), .Y(n3502) );
  OAI22XL U1934 ( .A0(n4056), .A1(n686), .B0(n1689), .B1(n4043), .Y(n3374) );
  OAI22XL U1935 ( .A0(n4060), .A1(n558), .B0(n1689), .B1(n4069), .Y(n3246) );
  OAI22XL U1936 ( .A0(n4079), .A1(n430), .B0(n1689), .B1(n4077), .Y(n3118) );
  OAI22XL U1937 ( .A0(n4094), .A1(n302), .B0(n1689), .B1(n4084), .Y(n2990) );
  OAI22XL U1938 ( .A0(n4108), .A1(n174), .B0(n1689), .B1(n4098), .Y(n2862) );
  OAI22XL U1939 ( .A0(n4186), .A1(n1070), .B0(n1689), .B1(n4177), .Y(n3758) );
  OAI22XL U1940 ( .A0(n4036), .A1(n797), .B0(n1672), .B1(n4029), .Y(n3485) );
  OAI22XL U1941 ( .A0(n4050), .A1(n669), .B0(n1672), .B1(n4044), .Y(n3357) );
  OAI22XL U1942 ( .A0(n4058), .A1(n541), .B0(n1672), .B1(n4069), .Y(n3229) );
  OAI22XL U1943 ( .A0(n4080), .A1(n413), .B0(n1672), .B1(n4076), .Y(n3101) );
  OAI22XL U1944 ( .A0(n4091), .A1(n285), .B0(n1672), .B1(n4085), .Y(n2973) );
  OAI22XL U1945 ( .A0(n4105), .A1(n157), .B0(n1672), .B1(n4099), .Y(n2845) );
  OAI22XL U1946 ( .A0(n4185), .A1(n1053), .B0(n1672), .B1(n4178), .Y(n3741) );
  OAI22XL U1947 ( .A0(n4037), .A1(n796), .B0(n1671), .B1(n4030), .Y(n3484) );
  OAI22XL U1948 ( .A0(n4051), .A1(n668), .B0(n1671), .B1(n4045), .Y(n3356) );
  OAI22XL U1949 ( .A0(n4057), .A1(n540), .B0(n1671), .B1(n4069), .Y(n3228) );
  OAI22XL U1950 ( .A0(n4080), .A1(n412), .B0(n1671), .B1(n4075), .Y(n3100) );
  OAI22XL U1951 ( .A0(n4092), .A1(n284), .B0(n1671), .B1(n4087), .Y(n2972) );
  OAI22XL U1952 ( .A0(n4106), .A1(n156), .B0(n1671), .B1(n4100), .Y(n2844) );
  OAI22XL U1953 ( .A0(n4185), .A1(n1052), .B0(n1671), .B1(n4178), .Y(n3740) );
  OAI22XL U1954 ( .A0(n4037), .A1(n795), .B0(n1670), .B1(n4030), .Y(n3483) );
  OAI22XL U1955 ( .A0(n4053), .A1(n667), .B0(n1670), .B1(n4045), .Y(n3355) );
  OAI22XL U1956 ( .A0(n4057), .A1(n539), .B0(n1670), .B1(n4069), .Y(n3227) );
  OAI22XL U1957 ( .A0(n4080), .A1(n411), .B0(n1670), .B1(n4076), .Y(n3099) );
  OAI22XL U1958 ( .A0(n4092), .A1(n283), .B0(n1670), .B1(n4087), .Y(n2971) );
  OAI22XL U1959 ( .A0(n4106), .A1(n155), .B0(n1670), .B1(n4100), .Y(n2843) );
  OAI22XL U1960 ( .A0(n4185), .A1(n1051), .B0(n1670), .B1(n4178), .Y(n3739) );
  OAI22XL U1961 ( .A0(n4037), .A1(n794), .B0(n1669), .B1(n4030), .Y(n3482) );
  OAI22XL U1962 ( .A0(n4055), .A1(n666), .B0(n1669), .B1(n4045), .Y(n3354) );
  OAI22XL U1963 ( .A0(n4057), .A1(n538), .B0(n1669), .B1(n4069), .Y(n3226) );
  OAI22XL U1964 ( .A0(n4080), .A1(n410), .B0(n1669), .B1(n4075), .Y(n3098) );
  OAI22XL U1965 ( .A0(n4092), .A1(n282), .B0(n1669), .B1(n4087), .Y(n2970) );
  OAI22XL U1966 ( .A0(n4106), .A1(n154), .B0(n1669), .B1(n4100), .Y(n2842) );
  OAI22XL U1967 ( .A0(n4185), .A1(n1050), .B0(n1669), .B1(n4178), .Y(n3738) );
  OAI22XL U1968 ( .A0(n4037), .A1(n793), .B0(n1668), .B1(n4030), .Y(n3481) );
  OAI22XL U1969 ( .A0(n4054), .A1(n665), .B0(n1668), .B1(n4045), .Y(n3353) );
  OAI22XL U1970 ( .A0(n4057), .A1(n537), .B0(n1668), .B1(n4069), .Y(n3225) );
  OAI22XL U1971 ( .A0(n4080), .A1(n409), .B0(n1668), .B1(n4076), .Y(n3097) );
  OAI22XL U1972 ( .A0(n4092), .A1(n281), .B0(n1668), .B1(n4087), .Y(n2969) );
  OAI22XL U1973 ( .A0(n4106), .A1(n153), .B0(n1668), .B1(n4100), .Y(n2841) );
  OAI22XL U1974 ( .A0(n4185), .A1(n1049), .B0(n1668), .B1(n4178), .Y(n3737) );
  OAI22XL U1975 ( .A0(n4037), .A1(n792), .B0(n1667), .B1(n4030), .Y(n3480) );
  OAI22XL U1976 ( .A0(n4056), .A1(n664), .B0(n1667), .B1(n4045), .Y(n3352) );
  OAI22XL U1977 ( .A0(n4058), .A1(n536), .B0(n1667), .B1(n4069), .Y(n3224) );
  OAI22XL U1978 ( .A0(n4080), .A1(n408), .B0(n1667), .B1(n4075), .Y(n3096) );
  OAI22XL U1979 ( .A0(n4092), .A1(n280), .B0(n1667), .B1(n4087), .Y(n2968) );
  OAI22XL U1980 ( .A0(n4106), .A1(n152), .B0(n1667), .B1(n4100), .Y(n2840) );
  OAI22XL U1981 ( .A0(n4185), .A1(n1048), .B0(n1667), .B1(n4178), .Y(n3736) );
  OAI22XL U1982 ( .A0(n4037), .A1(n791), .B0(n1666), .B1(n4030), .Y(n3479) );
  OAI22XL U1983 ( .A0(n4050), .A1(n663), .B0(n1666), .B1(n4045), .Y(n3351) );
  OAI22XL U1984 ( .A0(n4058), .A1(n535), .B0(n1666), .B1(n4069), .Y(n3223) );
  OAI22XL U1985 ( .A0(n4080), .A1(n407), .B0(n1666), .B1(n4076), .Y(n3095) );
  OAI22XL U1986 ( .A0(n4092), .A1(n279), .B0(n1666), .B1(n4087), .Y(n2967) );
  OAI22XL U1987 ( .A0(n4106), .A1(n151), .B0(n1666), .B1(n4100), .Y(n2839) );
  OAI22XL U1988 ( .A0(n4185), .A1(n1047), .B0(n1666), .B1(n4178), .Y(n3735) );
  OAI22XL U1989 ( .A0(n4037), .A1(n790), .B0(n1665), .B1(n4030), .Y(n3478) );
  OAI22XL U1990 ( .A0(n4051), .A1(n662), .B0(n1665), .B1(n4045), .Y(n3350) );
  OAI22XL U1991 ( .A0(n4058), .A1(n534), .B0(n1665), .B1(n4069), .Y(n3222) );
  OAI22XL U1992 ( .A0(n4081), .A1(n406), .B0(n1665), .B1(n4075), .Y(n3094) );
  OAI22XL U1993 ( .A0(n4092), .A1(n278), .B0(n1665), .B1(n4083), .Y(n2966) );
  OAI22XL U1994 ( .A0(n4106), .A1(n150), .B0(n1665), .B1(n4100), .Y(n2838) );
  OAI22XL U1995 ( .A0(n4186), .A1(n1046), .B0(n1665), .B1(n4179), .Y(n3734) );
  OAI22XL U1996 ( .A0(n4037), .A1(n789), .B0(n1664), .B1(n4030), .Y(n3477) );
  OAI22XL U1997 ( .A0(n4053), .A1(n661), .B0(n1664), .B1(n4045), .Y(n3349) );
  OAI22XL U1998 ( .A0(n4058), .A1(n533), .B0(n1664), .B1(n4068), .Y(n3221) );
  OAI22XL U1999 ( .A0(n4081), .A1(n405), .B0(n1664), .B1(n4073), .Y(n3093) );
  OAI22XL U2000 ( .A0(n4092), .A1(n277), .B0(n1664), .B1(n4087), .Y(n2965) );
  OAI22XL U2001 ( .A0(n4106), .A1(n149), .B0(n1664), .B1(n4100), .Y(n2837) );
  OAI22XL U2002 ( .A0(n4186), .A1(n1045), .B0(n1664), .B1(n4179), .Y(n3733) );
  OAI22XL U2003 ( .A0(n4037), .A1(n788), .B0(n1663), .B1(n4030), .Y(n3476) );
  OAI22XL U2004 ( .A0(n4055), .A1(n660), .B0(n1663), .B1(n4045), .Y(n3348) );
  OAI22XL U2005 ( .A0(n4058), .A1(n532), .B0(n1663), .B1(n4068), .Y(n3220) );
  OAI22XL U2006 ( .A0(n4081), .A1(n404), .B0(n1663), .B1(n4072), .Y(n3092) );
  OAI22XL U2007 ( .A0(n4092), .A1(n276), .B0(n1663), .B1(n4083), .Y(n2964) );
  OAI22XL U2008 ( .A0(n4106), .A1(n148), .B0(n1663), .B1(n4100), .Y(n2836) );
  OAI22XL U2009 ( .A0(n4186), .A1(n1044), .B0(n1663), .B1(n4179), .Y(n3732) );
  OAI22XL U2010 ( .A0(n4037), .A1(n787), .B0(n1662), .B1(n4030), .Y(n3475) );
  OAI22XL U2011 ( .A0(n4054), .A1(n659), .B0(n1662), .B1(n4045), .Y(n3347) );
  OAI22XL U2012 ( .A0(n4058), .A1(n531), .B0(n1662), .B1(n4068), .Y(n3219) );
  OAI22XL U2013 ( .A0(n4081), .A1(n403), .B0(n1662), .B1(n4075), .Y(n3091) );
  OAI22XL U2014 ( .A0(n4092), .A1(n275), .B0(n1662), .B1(n4089), .Y(n2963) );
  OAI22XL U2015 ( .A0(n4106), .A1(n147), .B0(n1662), .B1(n4100), .Y(n2835) );
  OAI22XL U2016 ( .A0(n4186), .A1(n1043), .B0(n1662), .B1(n4179), .Y(n3731) );
  OAI22XL U2017 ( .A0(n4037), .A1(n786), .B0(n1661), .B1(n4030), .Y(n3474) );
  OAI22XL U2018 ( .A0(n4050), .A1(n658), .B0(n1661), .B1(n4045), .Y(n3346) );
  OAI22XL U2019 ( .A0(n4058), .A1(n530), .B0(n1661), .B1(n4068), .Y(n3218) );
  OAI22XL U2020 ( .A0(n4081), .A1(n402), .B0(n1661), .B1(n4075), .Y(n3090) );
  OAI22XL U2021 ( .A0(n4092), .A1(n274), .B0(n1661), .B1(n4086), .Y(n2962) );
  OAI22XL U2022 ( .A0(n4106), .A1(n146), .B0(n1661), .B1(n4100), .Y(n2834) );
  OAI22XL U2023 ( .A0(n4186), .A1(n1042), .B0(n1661), .B1(n4179), .Y(n3730) );
  OAI22XL U2024 ( .A0(n4037), .A1(n785), .B0(n1660), .B1(n4030), .Y(n3473) );
  OAI22XL U2025 ( .A0(n4051), .A1(n657), .B0(n1660), .B1(n4045), .Y(n3345) );
  OAI22XL U2026 ( .A0(n4058), .A1(n529), .B0(n1660), .B1(n4068), .Y(n3217) );
  OAI22XL U2027 ( .A0(n4081), .A1(n401), .B0(n1660), .B1(n4075), .Y(n3089) );
  OAI22XL U2028 ( .A0(n4092), .A1(n273), .B0(n1660), .B1(n4083), .Y(n2961) );
  OAI22XL U2029 ( .A0(n4106), .A1(n145), .B0(n1660), .B1(n4100), .Y(n2833) );
  OAI22XL U2030 ( .A0(n4186), .A1(n1041), .B0(n1660), .B1(n4179), .Y(n3729) );
  OAI22XL U2031 ( .A0(n4038), .A1(n784), .B0(n1659), .B1(n4031), .Y(n3472) );
  OAI22XL U2032 ( .A0(n4052), .A1(n656), .B0(n1659), .B1(n4046), .Y(n3344) );
  OAI22XL U2033 ( .A0(n4058), .A1(n528), .B0(n1659), .B1(n4068), .Y(n3216) );
  OAI22XL U2034 ( .A0(n4081), .A1(n400), .B0(n1659), .B1(n4075), .Y(n3088) );
  OAI22XL U2035 ( .A0(n4093), .A1(n272), .B0(n1659), .B1(n4086), .Y(n2960) );
  OAI22XL U2036 ( .A0(n4107), .A1(n144), .B0(n1659), .B1(n4099), .Y(n2832) );
  OAI22XL U2037 ( .A0(n4186), .A1(n1040), .B0(n1659), .B1(n4179), .Y(n3728) );
  OAI22XL U2038 ( .A0(n4038), .A1(n783), .B0(n1658), .B1(n4031), .Y(n3471) );
  OAI22XL U2039 ( .A0(n4052), .A1(n655), .B0(n1658), .B1(n4046), .Y(n3343) );
  OAI22XL U2040 ( .A0(n4058), .A1(n527), .B0(n1658), .B1(n4068), .Y(n3215) );
  OAI22XL U2041 ( .A0(n4081), .A1(n399), .B0(n1658), .B1(n4075), .Y(n3087) );
  OAI22XL U2042 ( .A0(n4093), .A1(n271), .B0(n1658), .B1(n4086), .Y(n2959) );
  OAI22XL U2043 ( .A0(n4107), .A1(n143), .B0(n1658), .B1(n4097), .Y(n2831) );
  OAI22XL U2044 ( .A0(n4186), .A1(n1039), .B0(n1658), .B1(n4179), .Y(n3727) );
  OAI22XL U2045 ( .A0(n4038), .A1(n782), .B0(n1657), .B1(n4031), .Y(n3470) );
  OAI22XL U2046 ( .A0(n4052), .A1(n654), .B0(n1657), .B1(n4046), .Y(n3342) );
  OAI22XL U2047 ( .A0(n4058), .A1(n526), .B0(n1657), .B1(n4068), .Y(n3214) );
  OAI22XL U2048 ( .A0(n4081), .A1(n398), .B0(n1657), .B1(n4075), .Y(n3086) );
  OAI22XL U2049 ( .A0(n4093), .A1(n270), .B0(n1657), .B1(n4086), .Y(n2958) );
  OAI22XL U2050 ( .A0(n4107), .A1(n142), .B0(n1657), .B1(n4100), .Y(n2830) );
  OAI22XL U2051 ( .A0(n4186), .A1(n1038), .B0(n1657), .B1(n4179), .Y(n3726) );
  OAI22XL U2052 ( .A0(n4038), .A1(n781), .B0(n1656), .B1(n4031), .Y(n3469) );
  OAI22XL U2053 ( .A0(n4052), .A1(n653), .B0(n1656), .B1(n4046), .Y(n3341) );
  OAI22XL U2054 ( .A0(n4058), .A1(n525), .B0(n1656), .B1(n4068), .Y(n3213) );
  OAI22XL U2055 ( .A0(n4081), .A1(n397), .B0(n1656), .B1(n4075), .Y(n3085) );
  OAI22XL U2056 ( .A0(n4093), .A1(n269), .B0(n1656), .B1(n4086), .Y(n2957) );
  OAI22XL U2057 ( .A0(n4107), .A1(n141), .B0(n1656), .B1(n4101), .Y(n2829) );
  OAI22XL U2058 ( .A0(n4186), .A1(n1037), .B0(n1656), .B1(n4179), .Y(n3725) );
  OAI22XL U2059 ( .A0(n4038), .A1(n780), .B0(n1655), .B1(n4031), .Y(n3468) );
  OAI22XL U2060 ( .A0(n4053), .A1(n652), .B0(n1655), .B1(n4046), .Y(n3340) );
  OAI22XL U2061 ( .A0(n4059), .A1(n524), .B0(n1655), .B1(n4068), .Y(n3212) );
  OAI22XL U2062 ( .A0(n4081), .A1(n396), .B0(n1655), .B1(n4075), .Y(n3084) );
  OAI22XL U2063 ( .A0(n4093), .A1(n268), .B0(n1655), .B1(n4086), .Y(n2956) );
  OAI22XL U2064 ( .A0(n4107), .A1(n140), .B0(n1655), .B1(n4098), .Y(n2828) );
  OAI22XL U2065 ( .A0(n4186), .A1(n1036), .B0(n1655), .B1(n4179), .Y(n3724) );
  OAI22XL U2066 ( .A0(n4038), .A1(n779), .B0(n1654), .B1(n4031), .Y(n3467) );
  OAI22XL U2067 ( .A0(n4055), .A1(n651), .B0(n1654), .B1(n4046), .Y(n3339) );
  OAI22XL U2068 ( .A0(n4059), .A1(n523), .B0(n1654), .B1(n4068), .Y(n3211) );
  OAI22XL U2069 ( .A0(n4081), .A1(n395), .B0(n1654), .B1(n4075), .Y(n3083) );
  OAI22XL U2070 ( .A0(n4093), .A1(n267), .B0(n1654), .B1(n4086), .Y(n2955) );
  OAI22XL U2071 ( .A0(n4107), .A1(n139), .B0(n1654), .B1(n4097), .Y(n2827) );
  OAI22XL U2072 ( .A0(n4186), .A1(n1035), .B0(n1654), .B1(n4179), .Y(n3723) );
  OAI22XL U2073 ( .A0(n4038), .A1(n778), .B0(n1653), .B1(n4031), .Y(n3466) );
  OAI22XL U2074 ( .A0(n4051), .A1(n650), .B0(n1653), .B1(n4046), .Y(n3338) );
  OAI22XL U2075 ( .A0(n4059), .A1(n522), .B0(n1653), .B1(n4068), .Y(n3210) );
  OAI22XL U2076 ( .A0(n4082), .A1(n394), .B0(n1653), .B1(n4075), .Y(n3082) );
  OAI22XL U2077 ( .A0(n4093), .A1(n266), .B0(n1653), .B1(n4086), .Y(n2954) );
  OAI22XL U2078 ( .A0(n4107), .A1(n138), .B0(n1653), .B1(n4098), .Y(n2826) );
  OAI22XL U2079 ( .A0(n4187), .A1(n1034), .B0(n1653), .B1(n4180), .Y(n3722) );
  OAI22XL U2080 ( .A0(n4038), .A1(n777), .B0(n1652), .B1(n4031), .Y(n3465) );
  OAI22XL U2081 ( .A0(n4050), .A1(n649), .B0(n1652), .B1(n4046), .Y(n3337) );
  OAI22XL U2082 ( .A0(n4059), .A1(n521), .B0(n1652), .B1(n4068), .Y(n3209) );
  OAI22XL U2083 ( .A0(n4079), .A1(n393), .B0(n1652), .B1(n4075), .Y(n3081) );
  OAI22XL U2084 ( .A0(n4093), .A1(n265), .B0(n1652), .B1(n4086), .Y(n2953) );
  OAI22XL U2085 ( .A0(n4107), .A1(n137), .B0(n1652), .B1(n4097), .Y(n2825) );
  OAI22XL U2086 ( .A0(n4187), .A1(n1033), .B0(n1652), .B1(n4180), .Y(n3721) );
  OAI22XL U2087 ( .A0(n4038), .A1(n776), .B0(n1651), .B1(n4031), .Y(n3464) );
  OAI22XL U2088 ( .A0(n4054), .A1(n648), .B0(n1651), .B1(n4046), .Y(n3336) );
  OAI22XL U2089 ( .A0(n4059), .A1(n520), .B0(n1651), .B1(n4067), .Y(n3208) );
  OAI22XL U2090 ( .A0(n4078), .A1(n392), .B0(n1651), .B1(n4075), .Y(n3080) );
  OAI22XL U2091 ( .A0(n4093), .A1(n264), .B0(n1651), .B1(n4086), .Y(n2952) );
  OAI22XL U2092 ( .A0(n4107), .A1(n136), .B0(n1651), .B1(n4098), .Y(n2824) );
  OAI22XL U2093 ( .A0(n4187), .A1(n1032), .B0(n1651), .B1(n4180), .Y(n3720) );
  OAI22XL U2094 ( .A0(n4038), .A1(n775), .B0(n1650), .B1(n4031), .Y(n3463) );
  OAI22XL U2095 ( .A0(n4050), .A1(n647), .B0(n1650), .B1(n4046), .Y(n3335) );
  OAI22XL U2096 ( .A0(n4059), .A1(n519), .B0(n1650), .B1(n4067), .Y(n3207) );
  OAI22XL U2097 ( .A0(n4080), .A1(n391), .B0(n1650), .B1(n4075), .Y(n3079) );
  OAI22XL U2098 ( .A0(n4093), .A1(n263), .B0(n1650), .B1(n4086), .Y(n2951) );
  OAI22XL U2099 ( .A0(n4107), .A1(n135), .B0(n1650), .B1(n4097), .Y(n2823) );
  OAI22XL U2100 ( .A0(n4187), .A1(n1031), .B0(n1650), .B1(n4180), .Y(n3719) );
  OAI22XL U2101 ( .A0(n4038), .A1(n774), .B0(n1649), .B1(n4031), .Y(n3462) );
  OAI22XL U2102 ( .A0(n1700), .A1(n646), .B0(n1649), .B1(n4046), .Y(n3334) );
  OAI22XL U2103 ( .A0(n4059), .A1(n518), .B0(n1649), .B1(n4067), .Y(n3206) );
  OAI22XL U2104 ( .A0(n4079), .A1(n390), .B0(n1649), .B1(n4074), .Y(n3078) );
  OAI22XL U2105 ( .A0(n4093), .A1(n262), .B0(n1649), .B1(n4086), .Y(n2950) );
  OAI22XL U2106 ( .A0(n4107), .A1(n134), .B0(n1649), .B1(n4098), .Y(n2822) );
  OAI22XL U2107 ( .A0(n4187), .A1(n1030), .B0(n1649), .B1(n4180), .Y(n3718) );
  OAI22XL U2108 ( .A0(n4038), .A1(n773), .B0(n1648), .B1(n4031), .Y(n3461) );
  OAI22XL U2109 ( .A0(n4056), .A1(n645), .B0(n1648), .B1(n4046), .Y(n3333) );
  OAI22XL U2110 ( .A0(n4059), .A1(n517), .B0(n1648), .B1(n4067), .Y(n3205) );
  OAI22XL U2111 ( .A0(n4080), .A1(n389), .B0(n1648), .B1(n4074), .Y(n3077) );
  OAI22XL U2112 ( .A0(n4093), .A1(n261), .B0(n1648), .B1(n4086), .Y(n2949) );
  OAI22XL U2113 ( .A0(n4107), .A1(n133), .B0(n1648), .B1(n4097), .Y(n2821) );
  OAI22XL U2114 ( .A0(n4187), .A1(n1029), .B0(n1648), .B1(n4180), .Y(n3717) );
  OAI22XL U2115 ( .A0(n4039), .A1(n772), .B0(n1647), .B1(n4032), .Y(n3460) );
  OAI22XL U2116 ( .A0(n4051), .A1(n644), .B0(n1647), .B1(n4047), .Y(n3332) );
  OAI22XL U2117 ( .A0(n4059), .A1(n516), .B0(n1647), .B1(n4067), .Y(n3204) );
  OAI22XL U2118 ( .A0(n4081), .A1(n388), .B0(n1647), .B1(n4074), .Y(n3076) );
  OAI22XL U2119 ( .A0(n4091), .A1(n260), .B0(n1647), .B1(n4084), .Y(n2948) );
  OAI22XL U2120 ( .A0(n4105), .A1(n132), .B0(n1647), .B1(n4101), .Y(n2820) );
  OAI22XL U2121 ( .A0(n4187), .A1(n1028), .B0(n1647), .B1(n4180), .Y(n3716) );
  OAI22XL U2122 ( .A0(n4039), .A1(n771), .B0(n1646), .B1(n4032), .Y(n3459) );
  OAI22XL U2123 ( .A0(n4051), .A1(n643), .B0(n1646), .B1(n4047), .Y(n3331) );
  OAI22XL U2124 ( .A0(n4059), .A1(n515), .B0(n1646), .B1(n4067), .Y(n3203) );
  OAI22XL U2125 ( .A0(n4082), .A1(n387), .B0(n1646), .B1(n4074), .Y(n3075) );
  OAI22XL U2126 ( .A0(n4092), .A1(n259), .B0(n1646), .B1(n4084), .Y(n2947) );
  OAI22XL U2127 ( .A0(n4109), .A1(n131), .B0(n1646), .B1(n4101), .Y(n2819) );
  OAI22XL U2128 ( .A0(n4187), .A1(n1027), .B0(n1646), .B1(n4180), .Y(n3715) );
  OAI22XL U2129 ( .A0(n4039), .A1(n770), .B0(n1645), .B1(n4032), .Y(n3458) );
  OAI22XL U2130 ( .A0(n4051), .A1(n642), .B0(n1645), .B1(n4047), .Y(n3330) );
  OAI22XL U2131 ( .A0(n4059), .A1(n514), .B0(n1645), .B1(n4067), .Y(n3202) );
  OAI22XL U2132 ( .A0(n4079), .A1(n386), .B0(n1645), .B1(n4074), .Y(n3074) );
  OAI22XL U2133 ( .A0(n4095), .A1(n258), .B0(n1645), .B1(n4084), .Y(n2946) );
  OAI22XL U2134 ( .A0(n4105), .A1(n130), .B0(n1645), .B1(n4101), .Y(n2818) );
  OAI22XL U2135 ( .A0(n4187), .A1(n1026), .B0(n1645), .B1(n4180), .Y(n3714) );
  OAI22XL U2136 ( .A0(n4039), .A1(n769), .B0(n1644), .B1(n4032), .Y(n3457) );
  OAI22XL U2137 ( .A0(n4051), .A1(n641), .B0(n1644), .B1(n4047), .Y(n3329) );
  OAI22XL U2138 ( .A0(n4059), .A1(n513), .B0(n1644), .B1(n4067), .Y(n3201) );
  OAI22XL U2139 ( .A0(n4080), .A1(n385), .B0(n1644), .B1(n4074), .Y(n3073) );
  OAI22XL U2140 ( .A0(n4096), .A1(n257), .B0(n1644), .B1(n4084), .Y(n2945) );
  OAI22XL U2141 ( .A0(n4106), .A1(n129), .B0(n1644), .B1(n4101), .Y(n2817) );
  OAI22XL U2142 ( .A0(n4187), .A1(n1025), .B0(n1644), .B1(n4180), .Y(n3713) );
  OAI22XL U2143 ( .A0(n4039), .A1(n768), .B0(n1643), .B1(n4032), .Y(n3456) );
  OAI22XL U2144 ( .A0(n4051), .A1(n640), .B0(n1643), .B1(n4047), .Y(n3328) );
  OAI22XL U2145 ( .A0(n4060), .A1(n512), .B0(n1643), .B1(n4067), .Y(n3200) );
  OAI22XL U2146 ( .A0(n4081), .A1(n384), .B0(n1643), .B1(n4074), .Y(n3072) );
  OAI22XL U2147 ( .A0(n4094), .A1(n256), .B0(n1643), .B1(n4084), .Y(n2944) );
  OAI22XL U2148 ( .A0(n4110), .A1(n128), .B0(n1643), .B1(n4101), .Y(n2816) );
  OAI22XL U2149 ( .A0(n4187), .A1(n1024), .B0(n1643), .B1(n4180), .Y(n3712) );
  OAI22XL U2150 ( .A0(n4039), .A1(n767), .B0(n1642), .B1(n4032), .Y(n3455) );
  OAI22XL U2151 ( .A0(n4051), .A1(n639), .B0(n1642), .B1(n4047), .Y(n3327) );
  OAI22XL U2152 ( .A0(n4060), .A1(n511), .B0(n1642), .B1(n4067), .Y(n3199) );
  OAI22XL U2153 ( .A0(n4082), .A1(n383), .B0(n1642), .B1(n4074), .Y(n3071) );
  OAI22XL U2154 ( .A0(n4091), .A1(n255), .B0(n1642), .B1(n4084), .Y(n2943) );
  OAI22XL U2155 ( .A0(n4107), .A1(n127), .B0(n1642), .B1(n4101), .Y(n2815) );
  OAI22XL U2156 ( .A0(n4187), .A1(n1023), .B0(n1642), .B1(n4180), .Y(n3711) );
  OAI22XL U2157 ( .A0(n4039), .A1(n766), .B0(n1641), .B1(n4032), .Y(n3454) );
  OAI22XL U2158 ( .A0(n4051), .A1(n638), .B0(n1641), .B1(n4047), .Y(n3326) );
  OAI22XL U2159 ( .A0(n4060), .A1(n510), .B0(n1641), .B1(n4067), .Y(n3198) );
  OAI22XL U2160 ( .A0(n4080), .A1(n382), .B0(n1641), .B1(n4074), .Y(n3070) );
  OAI22XL U2161 ( .A0(n4090), .A1(n254), .B0(n1641), .B1(n4089), .Y(n2942) );
  OAI22XL U2162 ( .A0(n4108), .A1(n126), .B0(n1641), .B1(n4101), .Y(n2814) );
  OAI22XL U2163 ( .A0(n4188), .A1(n1022), .B0(n1641), .B1(n4183), .Y(n3710) );
  OAI22XL U2164 ( .A0(n4039), .A1(n765), .B0(n1640), .B1(n4032), .Y(n3453) );
  OAI22XL U2165 ( .A0(n4051), .A1(n637), .B0(n1640), .B1(n4047), .Y(n3325) );
  OAI22XL U2166 ( .A0(n4060), .A1(n509), .B0(n1640), .B1(n4067), .Y(n3197) );
  OAI22XL U2167 ( .A0(n4081), .A1(n381), .B0(n1640), .B1(n4074), .Y(n3069) );
  OAI22XL U2168 ( .A0(n4090), .A1(n253), .B0(n1640), .B1(n4086), .Y(n2941) );
  OAI22XL U2169 ( .A0(n4104), .A1(n125), .B0(n1640), .B1(n4101), .Y(n2813) );
  OAI22XL U2170 ( .A0(n4188), .A1(n1021), .B0(n1640), .B1(n4178), .Y(n3709) );
  OAI22XL U2171 ( .A0(n4039), .A1(n764), .B0(n1639), .B1(n4032), .Y(n3452) );
  OAI22XL U2172 ( .A0(n4051), .A1(n636), .B0(n1639), .B1(n4047), .Y(n3324) );
  OAI22XL U2173 ( .A0(n4060), .A1(n508), .B0(n1639), .B1(n4067), .Y(n3196) );
  OAI22XL U2174 ( .A0(n4081), .A1(n380), .B0(n1639), .B1(n4074), .Y(n3068) );
  OAI22XL U2175 ( .A0(n4090), .A1(n252), .B0(n1639), .B1(n4083), .Y(n2940) );
  OAI22XL U2176 ( .A0(n4109), .A1(n124), .B0(n1639), .B1(n4101), .Y(n2812) );
  OAI22XL U2177 ( .A0(n4188), .A1(n1020), .B0(n1639), .B1(n4177), .Y(n3708) );
  OAI22XL U2178 ( .A0(n4039), .A1(n763), .B0(n1638), .B1(n4032), .Y(n3451) );
  OAI22XL U2179 ( .A0(n4051), .A1(n635), .B0(n1638), .B1(n4047), .Y(n3323) );
  OAI22XL U2180 ( .A0(n4060), .A1(n507), .B0(n1638), .B1(n4066), .Y(n3195) );
  OAI22XL U2181 ( .A0(n4080), .A1(n379), .B0(n1638), .B1(n4074), .Y(n3067) );
  OAI22XL U2182 ( .A0(n4090), .A1(n251), .B0(n1638), .B1(n4084), .Y(n2939) );
  OAI22XL U2183 ( .A0(n4105), .A1(n123), .B0(n1638), .B1(n4101), .Y(n2811) );
  OAI22XL U2184 ( .A0(n4188), .A1(n1019), .B0(n1638), .B1(n4179), .Y(n3707) );
  OAI22XL U2185 ( .A0(n4039), .A1(n762), .B0(n1637), .B1(n4032), .Y(n3450) );
  OAI22XL U2186 ( .A0(n4051), .A1(n634), .B0(n1637), .B1(n4047), .Y(n3322) );
  OAI22XL U2187 ( .A0(n4060), .A1(n506), .B0(n1637), .B1(n4066), .Y(n3194) );
  OAI22XL U2188 ( .A0(n4081), .A1(n378), .B0(n1637), .B1(n4074), .Y(n3066) );
  OAI22XL U2189 ( .A0(n4090), .A1(n250), .B0(n1637), .B1(n4089), .Y(n2938) );
  OAI22XL U2190 ( .A0(n4106), .A1(n122), .B0(n1637), .B1(n4101), .Y(n2810) );
  OAI22XL U2191 ( .A0(n4188), .A1(n1018), .B0(n1637), .B1(n4180), .Y(n3706) );
  OAI22XL U2192 ( .A0(n4039), .A1(n761), .B0(n1636), .B1(n4032), .Y(n3449) );
  OAI22XL U2193 ( .A0(n4051), .A1(n633), .B0(n1636), .B1(n4047), .Y(n3321) );
  OAI22XL U2194 ( .A0(n4060), .A1(n505), .B0(n1636), .B1(n4066), .Y(n3193) );
  OAI22XL U2195 ( .A0(n4082), .A1(n377), .B0(n1636), .B1(n4074), .Y(n3065) );
  OAI22XL U2196 ( .A0(n4093), .A1(n249), .B0(n1636), .B1(n4086), .Y(n2937) );
  OAI22XL U2197 ( .A0(n4110), .A1(n121), .B0(n1636), .B1(n4101), .Y(n2809) );
  OAI22XL U2198 ( .A0(n4188), .A1(n1017), .B0(n1636), .B1(n4182), .Y(n3705) );
  OAI22XL U2199 ( .A0(n4040), .A1(n760), .B0(n1635), .B1(n4033), .Y(n3448) );
  OAI22XL U2200 ( .A0(n4052), .A1(n632), .B0(n1635), .B1(n4049), .Y(n3320) );
  OAI22XL U2201 ( .A0(n4060), .A1(n504), .B0(n1635), .B1(n4066), .Y(n3192) );
  OAI22XL U2202 ( .A0(n4078), .A1(n376), .B0(n1635), .B1(n4074), .Y(n3064) );
  OAI22XL U2203 ( .A0(n4090), .A1(n248), .B0(n1635), .B1(n4083), .Y(n2936) );
  OAI22XL U2204 ( .A0(n4108), .A1(n120), .B0(n1635), .B1(n4099), .Y(n2808) );
  OAI22XL U2205 ( .A0(n4188), .A1(n1016), .B0(n1635), .B1(n4181), .Y(n3704) );
  OAI22XL U2206 ( .A0(n4040), .A1(n759), .B0(n1634), .B1(n4033), .Y(n3447) );
  OAI22XL U2207 ( .A0(n4052), .A1(n631), .B0(n1634), .B1(n4049), .Y(n3319) );
  OAI22XL U2208 ( .A0(n4060), .A1(n503), .B0(n1634), .B1(n4066), .Y(n3191) );
  OAI22XL U2209 ( .A0(n4079), .A1(n375), .B0(n1634), .B1(n4074), .Y(n3063) );
  OAI22XL U2210 ( .A0(n4090), .A1(n247), .B0(n1634), .B1(n4086), .Y(n2935) );
  OAI22XL U2211 ( .A0(n4108), .A1(n119), .B0(n1634), .B1(n4101), .Y(n2807) );
  OAI22XL U2212 ( .A0(n4188), .A1(n1015), .B0(n1634), .B1(n2), .Y(n3703) );
  OAI22XL U2213 ( .A0(n4040), .A1(n758), .B0(n1633), .B1(n4033), .Y(n3446) );
  OAI22XL U2214 ( .A0(n4052), .A1(n630), .B0(n1633), .B1(n4049), .Y(n3318) );
  OAI22XL U2215 ( .A0(n4060), .A1(n502), .B0(n1633), .B1(n4066), .Y(n3190) );
  OAI22XL U2216 ( .A0(n4082), .A1(n374), .B0(n1633), .B1(n4074), .Y(n3062) );
  OAI22XL U2217 ( .A0(n4090), .A1(n246), .B0(n1633), .B1(n4089), .Y(n2934) );
  OAI22XL U2218 ( .A0(n4108), .A1(n118), .B0(n1633), .B1(n4099), .Y(n2806) );
  OAI22XL U2219 ( .A0(n4188), .A1(n1014), .B0(n1633), .B1(n4181), .Y(n3702) );
  OAI22XL U2220 ( .A0(n4040), .A1(n757), .B0(n1632), .B1(n4033), .Y(n3445) );
  OAI22XL U2221 ( .A0(n4052), .A1(n629), .B0(n1632), .B1(n4049), .Y(n3317) );
  OAI22XL U2222 ( .A0(n4060), .A1(n501), .B0(n1632), .B1(n4066), .Y(n3189) );
  OAI22XL U2223 ( .A0(n4078), .A1(n373), .B0(n1632), .B1(n4074), .Y(n3061) );
  OAI22XL U2224 ( .A0(n1692), .A1(n245), .B0(n1632), .B1(n4083), .Y(n2933) );
  OAI22XL U2225 ( .A0(n4108), .A1(n117), .B0(n1632), .B1(n4101), .Y(n2805) );
  OAI22XL U2226 ( .A0(n4188), .A1(n1013), .B0(n1632), .B1(n4181), .Y(n3701) );
  OAI22XL U2227 ( .A0(n4040), .A1(n756), .B0(n1631), .B1(n4033), .Y(n3444) );
  OAI22XL U2228 ( .A0(n4052), .A1(n628), .B0(n1631), .B1(n4049), .Y(n3316) );
  OAI22XL U2229 ( .A0(n4062), .A1(n500), .B0(n1631), .B1(n4066), .Y(n3188) );
  OAI22XL U2230 ( .A0(n4078), .A1(n372), .B0(n1631), .B1(n4073), .Y(n3060) );
  OAI22XL U2231 ( .A0(n1692), .A1(n244), .B0(n1631), .B1(n4086), .Y(n2932) );
  OAI22XL U2232 ( .A0(n4108), .A1(n116), .B0(n1631), .B1(n4100), .Y(n2804) );
  OAI22XL U2233 ( .A0(n4188), .A1(n1012), .B0(n1631), .B1(n4181), .Y(n3700) );
  OAI22XL U2234 ( .A0(n4040), .A1(n755), .B0(n1630), .B1(n4033), .Y(n3443) );
  OAI22XL U2235 ( .A0(n4052), .A1(n627), .B0(n1630), .B1(n4049), .Y(n3315) );
  OAI22XL U2236 ( .A0(n4058), .A1(n499), .B0(n1630), .B1(n4066), .Y(n3187) );
  OAI22XL U2237 ( .A0(n4078), .A1(n371), .B0(n1630), .B1(n4072), .Y(n3059) );
  OAI22XL U2238 ( .A0(n1692), .A1(n243), .B0(n1630), .B1(n4089), .Y(n2931) );
  OAI22XL U2239 ( .A0(n4108), .A1(n115), .B0(n1630), .B1(n4097), .Y(n2803) );
  OAI22XL U2240 ( .A0(n4188), .A1(n1011), .B0(n1630), .B1(n4181), .Y(n3699) );
  OAI22XL U2241 ( .A0(n4040), .A1(n754), .B0(n1629), .B1(n4033), .Y(n3442) );
  OAI22XL U2242 ( .A0(n4052), .A1(n626), .B0(n1629), .B1(n4049), .Y(n3314) );
  OAI22XL U2243 ( .A0(n4059), .A1(n498), .B0(n1629), .B1(n4066), .Y(n3186) );
  OAI22XL U2244 ( .A0(n4080), .A1(n370), .B0(n1629), .B1(n4071), .Y(n3058) );
  OAI22XL U2245 ( .A0(n1692), .A1(n242), .B0(n1629), .B1(n4083), .Y(n2930) );
  OAI22XL U2246 ( .A0(n4108), .A1(n114), .B0(n1629), .B1(n4102), .Y(n2802) );
  OAI22XL U2247 ( .A0(n4188), .A1(n1010), .B0(n1629), .B1(n4179), .Y(n3698) );
  OAI22XL U2248 ( .A0(n4040), .A1(n753), .B0(n1628), .B1(n4033), .Y(n3441) );
  OAI22XL U2249 ( .A0(n4052), .A1(n625), .B0(n1628), .B1(n4049), .Y(n3313) );
  OAI22XL U2250 ( .A0(n4061), .A1(n497), .B0(n1628), .B1(n4066), .Y(n3185) );
  OAI22XL U2251 ( .A0(n4081), .A1(n369), .B0(n1628), .B1(n4077), .Y(n3057) );
  OAI22XL U2252 ( .A0(n1692), .A1(n241), .B0(n1628), .B1(n4086), .Y(n2929) );
  OAI22XL U2253 ( .A0(n4108), .A1(n113), .B0(n1628), .B1(n4098), .Y(n2801) );
  OAI22XL U2254 ( .A0(n4187), .A1(n1009), .B0(n1628), .B1(n4183), .Y(n3697) );
  OAI22XL U2255 ( .A0(n4040), .A1(n752), .B0(n1627), .B1(n4033), .Y(n3440) );
  OAI22XL U2256 ( .A0(n4052), .A1(n624), .B0(n1627), .B1(n4049), .Y(n3312) );
  OAI22XL U2257 ( .A0(n4060), .A1(n496), .B0(n1627), .B1(n4066), .Y(n3184) );
  OAI22XL U2258 ( .A0(n4081), .A1(n368), .B0(n1627), .B1(n4071), .Y(n3056) );
  OAI22XL U2259 ( .A0(n4090), .A1(n240), .B0(n1627), .B1(n4089), .Y(n2928) );
  OAI22XL U2260 ( .A0(n4108), .A1(n112), .B0(n1627), .B1(n4102), .Y(n2800) );
  OAI22XL U2261 ( .A0(n4188), .A1(n1008), .B0(n1627), .B1(n4177), .Y(n3696) );
  OAI22XL U2262 ( .A0(n4040), .A1(n751), .B0(n1626), .B1(n4033), .Y(n3439) );
  OAI22XL U2263 ( .A0(n4052), .A1(n623), .B0(n1626), .B1(n4049), .Y(n3311) );
  OAI22XL U2264 ( .A0(n4062), .A1(n495), .B0(n1626), .B1(n4065), .Y(n3183) );
  OAI22XL U2265 ( .A0(n4082), .A1(n367), .B0(n1626), .B1(n4075), .Y(n3055) );
  OAI22XL U2266 ( .A0(n4090), .A1(n239), .B0(n1626), .B1(n4083), .Y(n2927) );
  OAI22XL U2267 ( .A0(n4108), .A1(n111), .B0(n1626), .B1(n4097), .Y(n2799) );
  OAI22XL U2268 ( .A0(n4185), .A1(n1007), .B0(n1626), .B1(n4178), .Y(n3695) );
  OAI22XL U2269 ( .A0(n4040), .A1(n750), .B0(n1625), .B1(n4033), .Y(n3438) );
  OAI22XL U2270 ( .A0(n4052), .A1(n622), .B0(n1625), .B1(n4046), .Y(n3310) );
  OAI22XL U2271 ( .A0(n4058), .A1(n494), .B0(n1625), .B1(n4065), .Y(n3182) );
  OAI22XL U2272 ( .A0(n4079), .A1(n366), .B0(n1625), .B1(n4071), .Y(n3054) );
  OAI22XL U2273 ( .A0(n4090), .A1(n238), .B0(n1625), .B1(n4086), .Y(n2926) );
  OAI22XL U2274 ( .A0(n4108), .A1(n110), .B0(n1625), .B1(n4103), .Y(n2798) );
  OAI22XL U2275 ( .A0(n4186), .A1(n1006), .B0(n1625), .B1(n4179), .Y(n3694) );
  OAI22XL U2276 ( .A0(n4040), .A1(n749), .B0(n1624), .B1(n4033), .Y(n3437) );
  OAI22XL U2277 ( .A0(n4052), .A1(n621), .B0(n1624), .B1(n4043), .Y(n3309) );
  OAI22XL U2278 ( .A0(n4059), .A1(n493), .B0(n1624), .B1(n4065), .Y(n3181) );
  OAI22XL U2279 ( .A0(n4078), .A1(n365), .B0(n1624), .B1(n4072), .Y(n3053) );
  OAI22XL U2280 ( .A0(n4090), .A1(n237), .B0(n1624), .B1(n4089), .Y(n2925) );
  OAI22XL U2281 ( .A0(n4108), .A1(n109), .B0(n1624), .B1(n5), .Y(n2797) );
  OAI22XL U2282 ( .A0(n4189), .A1(n1005), .B0(n1624), .B1(n4183), .Y(n3693) );
  OAI22XL U2283 ( .A0(n4038), .A1(n748), .B0(n1623), .B1(n4030), .Y(n3436) );
  OAI22XL U2284 ( .A0(n4053), .A1(n620), .B0(n1623), .B1(n4048), .Y(n3308) );
  OAI22XL U2285 ( .A0(n4061), .A1(n492), .B0(n1623), .B1(n4065), .Y(n3180) );
  OAI22XL U2286 ( .A0(n4081), .A1(n364), .B0(n1623), .B1(n4077), .Y(n3052) );
  OAI22XL U2287 ( .A0(n4092), .A1(n236), .B0(n1623), .B1(n4087), .Y(n2924) );
  OAI22XL U2288 ( .A0(n4104), .A1(n108), .B0(n1623), .B1(n4103), .Y(n2796) );
  OAI22XL U2289 ( .A0(n4184), .A1(n1004), .B0(n1623), .B1(n4177), .Y(n3692) );
  OAI22XL U2290 ( .A0(n4036), .A1(n747), .B0(n1622), .B1(n4032), .Y(n3435) );
  OAI22XL U2291 ( .A0(n4053), .A1(n619), .B0(n1622), .B1(n4045), .Y(n3307) );
  OAI22XL U2292 ( .A0(n4061), .A1(n491), .B0(n1622), .B1(n4065), .Y(n3179) );
  OAI22XL U2293 ( .A0(n1694), .A1(n363), .B0(n1622), .B1(n4073), .Y(n3051) );
  OAI22XL U2294 ( .A0(n4095), .A1(n235), .B0(n1622), .B1(n4087), .Y(n2923) );
  OAI22XL U2295 ( .A0(n4106), .A1(n107), .B0(n1622), .B1(n4102), .Y(n2795) );
  OAI22XL U2296 ( .A0(n4189), .A1(n1003), .B0(n1622), .B1(n4178), .Y(n3691) );
  OAI22XL U2297 ( .A0(n4040), .A1(n746), .B0(n1621), .B1(n4033), .Y(n3434) );
  OAI22XL U2298 ( .A0(n4053), .A1(n618), .B0(n1621), .B1(n4047), .Y(n3306) );
  OAI22XL U2299 ( .A0(n4057), .A1(n490), .B0(n1621), .B1(n4065), .Y(n3178) );
  OAI22XL U2300 ( .A0(n4078), .A1(n362), .B0(n1621), .B1(n4072), .Y(n3050) );
  OAI22XL U2301 ( .A0(n4096), .A1(n234), .B0(n1621), .B1(n4087), .Y(n2922) );
  OAI22XL U2302 ( .A0(n4110), .A1(n106), .B0(n1621), .B1(n4103), .Y(n2794) );
  OAI22XL U2303 ( .A0(n4190), .A1(n1002), .B0(n1621), .B1(n4179), .Y(n3690) );
  OAI22XL U2304 ( .A0(n4042), .A1(n745), .B0(n1620), .B1(n4034), .Y(n3433) );
  OAI22XL U2305 ( .A0(n4053), .A1(n617), .B0(n1620), .B1(n4046), .Y(n3305) );
  OAI22XL U2306 ( .A0(n4057), .A1(n489), .B0(n1620), .B1(n4065), .Y(n3177) );
  OAI22XL U2307 ( .A0(n4078), .A1(n361), .B0(n1620), .B1(n4077), .Y(n3049) );
  OAI22XL U2308 ( .A0(n4096), .A1(n233), .B0(n1620), .B1(n4087), .Y(n2921) );
  OAI22XL U2309 ( .A0(n4107), .A1(n105), .B0(n1620), .B1(n4102), .Y(n2793) );
  OAI22XL U2310 ( .A0(n4187), .A1(n1001), .B0(n1620), .B1(n4183), .Y(n3689) );
  OAI22XL U2311 ( .A0(n4042), .A1(n744), .B0(n1619), .B1(n4031), .Y(n3432) );
  OAI22XL U2312 ( .A0(n4053), .A1(n616), .B0(n1619), .B1(n4043), .Y(n3304) );
  OAI22XL U2313 ( .A0(n4061), .A1(n488), .B0(n1619), .B1(n4065), .Y(n3176) );
  OAI22XL U2314 ( .A0(n4079), .A1(n360), .B0(n1619), .B1(n4073), .Y(n3048) );
  OAI22XL U2315 ( .A0(n4094), .A1(n232), .B0(n1619), .B1(n4087), .Y(n2920) );
  OAI22XL U2316 ( .A0(n4108), .A1(n104), .B0(n1619), .B1(n4103), .Y(n2792) );
  OAI22XL U2317 ( .A0(n4188), .A1(n1000), .B0(n1619), .B1(n4177), .Y(n3688) );
  OAI22XL U2318 ( .A0(n4038), .A1(n826), .B0(n1539), .B1(n4030), .Y(n3514) );
  OAI22XL U2319 ( .A0(n4052), .A1(n698), .B0(n1539), .B1(n4048), .Y(n3386) );
  OAI22XL U2320 ( .A0(n4060), .A1(n570), .B0(n1539), .B1(n4070), .Y(n3258) );
  OAI22XL U2321 ( .A0(n1694), .A1(n442), .B0(n1539), .B1(n4072), .Y(n3130) );
  OAI22XL U2322 ( .A0(n4090), .A1(n314), .B0(n1539), .B1(n4083), .Y(n3002) );
  OAI22XL U2323 ( .A0(n4109), .A1(n186), .B0(n1539), .B1(n4097), .Y(n2874) );
  OAI22XL U2324 ( .A0(n4189), .A1(n1082), .B0(n1539), .B1(n4183), .Y(n3770) );
  OAI22XL U2325 ( .A0(n4036), .A1(n825), .B0(n1538), .B1(n4032), .Y(n3513) );
  OAI22XL U2326 ( .A0(n4054), .A1(n697), .B0(n1538), .B1(n4047), .Y(n3385) );
  OAI22XL U2327 ( .A0(n4058), .A1(n569), .B0(n1538), .B1(n4070), .Y(n3257) );
  OAI22XL U2328 ( .A0(n4079), .A1(n441), .B0(n1538), .B1(n4077), .Y(n3129) );
  OAI22XL U2329 ( .A0(n4093), .A1(n313), .B0(n1538), .B1(n4083), .Y(n3001) );
  OAI22XL U2330 ( .A0(n4105), .A1(n185), .B0(n1538), .B1(n4097), .Y(n2873) );
  OAI22XL U2331 ( .A0(n4190), .A1(n1081), .B0(n1538), .B1(n4183), .Y(n3769) );
  OAI22XL U2332 ( .A0(n4036), .A1(n824), .B0(n1537), .B1(n4033), .Y(n3512) );
  OAI22XL U2333 ( .A0(n4056), .A1(n696), .B0(n1537), .B1(n4049), .Y(n3384) );
  OAI22XL U2334 ( .A0(n4059), .A1(n568), .B0(n1537), .B1(n4070), .Y(n3256) );
  OAI22XL U2335 ( .A0(n4079), .A1(n440), .B0(n1537), .B1(n4077), .Y(n3128) );
  OAI22XL U2336 ( .A0(n4093), .A1(n312), .B0(n1537), .B1(n4083), .Y(n3000) );
  OAI22XL U2337 ( .A0(n4104), .A1(n184), .B0(n1537), .B1(n4097), .Y(n2872) );
  OAI22XL U2338 ( .A0(n4187), .A1(n1080), .B0(n1537), .B1(n4183), .Y(n3768) );
  OAI22XL U2339 ( .A0(n4040), .A1(n823), .B0(n1536), .B1(n4035), .Y(n3511) );
  OAI22XL U2340 ( .A0(n4056), .A1(n695), .B0(n1536), .B1(n4), .Y(n3383) );
  OAI22XL U2341 ( .A0(n4062), .A1(n567), .B0(n1536), .B1(n4070), .Y(n3255) );
  OAI22XL U2342 ( .A0(n4082), .A1(n439), .B0(n1536), .B1(n4077), .Y(n3127) );
  OAI22XL U2343 ( .A0(n4090), .A1(n311), .B0(n1536), .B1(n4083), .Y(n2999) );
  OAI22XL U2344 ( .A0(n4104), .A1(n183), .B0(n1536), .B1(n4097), .Y(n2871) );
  OAI22XL U2345 ( .A0(n4188), .A1(n1079), .B0(n1536), .B1(n4183), .Y(n3767) );
  OAI22XL U2346 ( .A0(n1702), .A1(n822), .B0(n1535), .B1(n3), .Y(n3510) );
  OAI22XL U2347 ( .A0(n4052), .A1(n694), .B0(n1535), .B1(n4049), .Y(n3382) );
  OAI22XL U2348 ( .A0(n4061), .A1(n566), .B0(n1535), .B1(n4070), .Y(n3254) );
  OAI22XL U2349 ( .A0(n4082), .A1(n438), .B0(n1535), .B1(n4077), .Y(n3126) );
  OAI22XL U2350 ( .A0(n4093), .A1(n310), .B0(n1535), .B1(n4083), .Y(n2998) );
  OAI22XL U2351 ( .A0(n4104), .A1(n182), .B0(n1535), .B1(n4097), .Y(n2870) );
  OAI22XL U2352 ( .A0(n4187), .A1(n1078), .B0(n1535), .B1(n4177), .Y(n3766) );
  OAI22XL U2353 ( .A0(n4042), .A1(n821), .B0(n1534), .B1(n4035), .Y(n3509) );
  OAI22XL U2354 ( .A0(n4051), .A1(n693), .B0(n1534), .B1(n4049), .Y(n3381) );
  OAI22XL U2355 ( .A0(n4060), .A1(n565), .B0(n1534), .B1(n4070), .Y(n3253) );
  OAI22XL U2356 ( .A0(n4079), .A1(n437), .B0(n1534), .B1(n4077), .Y(n3125) );
  OAI22XL U2357 ( .A0(n4093), .A1(n309), .B0(n1534), .B1(n4083), .Y(n2997) );
  OAI22XL U2358 ( .A0(n4104), .A1(n181), .B0(n1534), .B1(n4097), .Y(n2869) );
  OAI22XL U2359 ( .A0(n4186), .A1(n1077), .B0(n1534), .B1(n4183), .Y(n3765) );
  OAI22XL U2360 ( .A0(n4038), .A1(n820), .B0(n1533), .B1(n4029), .Y(n3508) );
  OAI22XL U2361 ( .A0(n4056), .A1(n692), .B0(n1533), .B1(n4043), .Y(n3380) );
  OAI22XL U2362 ( .A0(n1699), .A1(n564), .B0(n1533), .B1(n4070), .Y(n3252) );
  OAI22XL U2363 ( .A0(n4082), .A1(n436), .B0(n1533), .B1(n4077), .Y(n3124) );
  OAI22XL U2364 ( .A0(n4091), .A1(n308), .B0(n1533), .B1(n4084), .Y(n2996) );
  OAI22XL U2365 ( .A0(n4109), .A1(n180), .B0(n1533), .B1(n4098), .Y(n2868) );
  OAI22XL U2366 ( .A0(n4185), .A1(n1076), .B0(n1533), .B1(n4179), .Y(n3764) );
  OAI22XL U2367 ( .A0(n4042), .A1(n819), .B0(n1532), .B1(n4029), .Y(n3507) );
  OAI22XL U2368 ( .A0(n4056), .A1(n691), .B0(n1532), .B1(n4043), .Y(n3379) );
  OAI22XL U2369 ( .A0(n1699), .A1(n563), .B0(n1532), .B1(n4070), .Y(n3251) );
  OAI22XL U2370 ( .A0(n4078), .A1(n435), .B0(n1532), .B1(n4077), .Y(n3123) );
  OAI22XL U2371 ( .A0(n4092), .A1(n307), .B0(n1532), .B1(n4084), .Y(n2995) );
  OAI22XL U2372 ( .A0(n4105), .A1(n179), .B0(n1532), .B1(n4098), .Y(n2867) );
  OAI22XL U2373 ( .A0(n4186), .A1(n1075), .B0(n1532), .B1(n4179), .Y(n3763) );
  OAI22XL U2374 ( .A0(n4042), .A1(n818), .B0(n1531), .B1(n4029), .Y(n3506) );
  OAI22XL U2375 ( .A0(n4056), .A1(n690), .B0(n1531), .B1(n4043), .Y(n3378) );
  OAI22XL U2376 ( .A0(n1699), .A1(n562), .B0(n1531), .B1(n4069), .Y(n3250) );
  OAI22XL U2377 ( .A0(n4078), .A1(n434), .B0(n1531), .B1(n4077), .Y(n3122) );
  OAI22XL U2378 ( .A0(n4095), .A1(n306), .B0(n1531), .B1(n4084), .Y(n2994) );
  OAI22XL U2379 ( .A0(n1578), .A1(n178), .B0(n1531), .B1(n4098), .Y(n2866) );
  OAI22XL U2380 ( .A0(n4189), .A1(n1074), .B0(n1531), .B1(n4179), .Y(n3762) );
  OAI22XL U2381 ( .A0(n4042), .A1(n817), .B0(n1530), .B1(n4029), .Y(n3505) );
  OAI22XL U2382 ( .A0(n1700), .A1(n689), .B0(n1530), .B1(n4043), .Y(n3377) );
  OAI22XL U2383 ( .A0(n1699), .A1(n561), .B0(n1530), .B1(n4069), .Y(n3249) );
  OAI22XL U2384 ( .A0(n4078), .A1(n433), .B0(n1530), .B1(n4077), .Y(n3121) );
  OAI22XL U2385 ( .A0(n4096), .A1(n305), .B0(n1530), .B1(n4084), .Y(n2993) );
  OAI22XL U2386 ( .A0(n4104), .A1(n177), .B0(n1530), .B1(n4098), .Y(n2865) );
  OAI22XL U2387 ( .A0(n4190), .A1(n1073), .B0(n1530), .B1(n4179), .Y(n3761) );
  OAI22XL U2388 ( .A0(n4042), .A1(n816), .B0(n1529), .B1(n4029), .Y(n3504) );
  OAI22XL U2389 ( .A0(n1700), .A1(n688), .B0(n1529), .B1(n4043), .Y(n3376) );
  OAI22XL U2390 ( .A0(n1699), .A1(n560), .B0(n1529), .B1(n4069), .Y(n3248) );
  OAI22XL U2391 ( .A0(n4078), .A1(n432), .B0(n1529), .B1(n4077), .Y(n3120) );
  OAI22XL U2392 ( .A0(n4095), .A1(n304), .B0(n1529), .B1(n4084), .Y(n2992) );
  OAI22XL U2393 ( .A0(n4104), .A1(n176), .B0(n1529), .B1(n4098), .Y(n2864) );
  OAI22XL U2394 ( .A0(n4184), .A1(n1072), .B0(n1529), .B1(n4178), .Y(n3760) );
  OAI22XL U2395 ( .A0(n1702), .A1(n815), .B0(n1527), .B1(n4029), .Y(n3503) );
  OAI22XL U2396 ( .A0(n1700), .A1(n687), .B0(n1527), .B1(n4043), .Y(n3375) );
  OAI22XL U2397 ( .A0(n4057), .A1(n559), .B0(n1527), .B1(n4069), .Y(n3247) );
  OAI22XL U2398 ( .A0(n1694), .A1(n431), .B0(n1527), .B1(n4077), .Y(n3119) );
  OAI22XL U2399 ( .A0(n4094), .A1(n303), .B0(n1527), .B1(n4084), .Y(n2991) );
  OAI22XL U2400 ( .A0(n4104), .A1(n175), .B0(n1527), .B1(n4098), .Y(n2863) );
  OAI22XL U2401 ( .A0(n4188), .A1(n1071), .B0(n1527), .B1(n4179), .Y(n3759) );
  OAI22XL U2402 ( .A0(n1611), .A1(n4028), .B0(n4018), .B1(n864), .Y(n3552) );
  OAI22XL U2403 ( .A0(n1611), .A1(n4072), .B0(n1339), .B1(n352), .Y(n3040) );
  OAI22XL U2404 ( .A0(n1610), .A1(n4028), .B0(n4019), .B1(n863), .Y(n3551) );
  OAI22XL U2405 ( .A0(n1610), .A1(n4072), .B0(n1338), .B1(n351), .Y(n3039) );
  OAI22XL U2406 ( .A0(n1609), .A1(n4028), .B0(n4020), .B1(n862), .Y(n3550) );
  OAI22XL U2407 ( .A0(n1609), .A1(n4072), .B0(n1339), .B1(n350), .Y(n3038) );
  OAI22XL U2408 ( .A0(n1608), .A1(n4028), .B0(n4020), .B1(n861), .Y(n3549) );
  OAI22XL U2409 ( .A0(n1608), .A1(n4072), .B0(n1338), .B1(n349), .Y(n3037) );
  OAI22XL U2410 ( .A0(n1607), .A1(n4028), .B0(n4021), .B1(n860), .Y(n3548) );
  OAI22XL U2411 ( .A0(n1607), .A1(n4072), .B0(n1339), .B1(n348), .Y(n3036) );
  OAI22XL U2412 ( .A0(n1606), .A1(n4028), .B0(n4021), .B1(n859), .Y(n3547) );
  OAI22XL U2413 ( .A0(n1606), .A1(n4076), .B0(n1338), .B1(n347), .Y(n3035) );
  OAI22XL U2414 ( .A0(n1605), .A1(n4028), .B0(n4021), .B1(n858), .Y(n3546) );
  OAI22XL U2415 ( .A0(n1605), .A1(n4076), .B0(n1339), .B1(n346), .Y(n3034) );
  OAI22XL U2416 ( .A0(n1604), .A1(n4028), .B0(n4021), .B1(n857), .Y(n3545) );
  OAI22XL U2417 ( .A0(n1604), .A1(n4077), .B0(n1338), .B1(n345), .Y(n3033) );
  OAI22XL U2418 ( .A0(n1603), .A1(n4028), .B0(n4021), .B1(n856), .Y(n3544) );
  OAI22XL U2419 ( .A0(n1603), .A1(n4072), .B0(n1339), .B1(n344), .Y(n3032) );
  OAI22XL U2420 ( .A0(n1589), .A1(n4028), .B0(n4016), .B1(n842), .Y(n3530) );
  OAI22XL U2421 ( .A0(n1589), .A1(n4064), .B0(n1698), .B1(n458), .Y(n3146) );
  OAI22XL U2422 ( .A0(n1588), .A1(n4023), .B0(n4016), .B1(n841), .Y(n3529) );
  OAI22XL U2423 ( .A0(n1588), .A1(n4064), .B0(n1698), .B1(n457), .Y(n3145) );
  OAI22XL U2424 ( .A0(n1587), .A1(n4024), .B0(n1706), .B1(n840), .Y(n3528) );
  OAI22XL U2425 ( .A0(n1587), .A1(n4064), .B0(n1698), .B1(n456), .Y(n3144) );
  OAI22XL U2426 ( .A0(n1586), .A1(n4025), .B0(n1706), .B1(n839), .Y(n3527) );
  OAI22XL U2427 ( .A0(n1586), .A1(n4064), .B0(n1698), .B1(n455), .Y(n3143) );
  OAI22XL U2428 ( .A0(n1585), .A1(n4024), .B0(n4021), .B1(n838), .Y(n3526) );
  OAI22XL U2429 ( .A0(n1585), .A1(n4064), .B0(n1698), .B1(n454), .Y(n3142) );
  OAI22XL U2430 ( .A0(n1584), .A1(n4025), .B0(n4021), .B1(n837), .Y(n3525) );
  OAI22XL U2431 ( .A0(n1584), .A1(n4064), .B0(n1698), .B1(n453), .Y(n3141) );
  OAI22XL U2432 ( .A0(n1583), .A1(n4026), .B0(n4021), .B1(n836), .Y(n3524) );
  OAI22XL U2433 ( .A0(n1583), .A1(n4064), .B0(n1698), .B1(n452), .Y(n3140) );
  OAI22XL U2434 ( .A0(n1582), .A1(n4023), .B0(n4021), .B1(n835), .Y(n3523) );
  OAI22XL U2435 ( .A0(n1582), .A1(n4064), .B0(n1698), .B1(n451), .Y(n3139) );
  OAI22XL U2436 ( .A0(n1581), .A1(n4022), .B0(n4021), .B1(n834), .Y(n3522) );
  OAI22XL U2437 ( .A0(n1581), .A1(n4064), .B0(n4063), .B1(n450), .Y(n3138) );
  OAI22XL U2438 ( .A0(n1579), .A1(n4028), .B0(n4021), .B1(n833), .Y(n3521) );
  OAI22XL U2439 ( .A0(n1579), .A1(n4066), .B0(n4063), .B1(n449), .Y(n3137) );
  OAI22XL U2440 ( .A0(n1688), .A1(n4022), .B0(n4016), .B1(n941), .Y(n3629) );
  OAI22XL U2441 ( .A0(n1688), .A1(n4064), .B0(n4063), .B1(n557), .Y(n3245) );
  OAI22XL U2442 ( .A0(n1687), .A1(n4022), .B0(n4016), .B1(n940), .Y(n3628) );
  OAI22XL U2443 ( .A0(n1687), .A1(n4068), .B0(n4063), .B1(n556), .Y(n3244) );
  OAI22XL U2444 ( .A0(n1686), .A1(n4022), .B0(n4016), .B1(n939), .Y(n3627) );
  OAI22XL U2445 ( .A0(n1686), .A1(n4067), .B0(n4063), .B1(n555), .Y(n3243) );
  OAI22XL U2446 ( .A0(n1685), .A1(n4022), .B0(n4016), .B1(n938), .Y(n3626) );
  OAI22XL U2447 ( .A0(n1685), .A1(n4065), .B0(n4063), .B1(n554), .Y(n3242) );
  OAI22XL U2448 ( .A0(n1684), .A1(n4022), .B0(n4017), .B1(n937), .Y(n3625) );
  OAI22XL U2449 ( .A0(n1684), .A1(n4064), .B0(n4063), .B1(n553), .Y(n3241) );
  OAI22XL U2450 ( .A0(n1683), .A1(n4023), .B0(n4017), .B1(n936), .Y(n3624) );
  OAI22XL U2451 ( .A0(n1683), .A1(n4068), .B0(n4063), .B1(n552), .Y(n3240) );
  OAI22XL U2452 ( .A0(n1682), .A1(n4023), .B0(n4017), .B1(n935), .Y(n3623) );
  OAI22XL U2453 ( .A0(n1682), .A1(n4067), .B0(n4063), .B1(n551), .Y(n3239) );
  OAI22XL U2454 ( .A0(n1681), .A1(n4023), .B0(n4017), .B1(n934), .Y(n3622) );
  OAI22XL U2455 ( .A0(n1681), .A1(n4066), .B0(n4063), .B1(n550), .Y(n3238) );
  OAI22XL U2456 ( .A0(n1680), .A1(n4023), .B0(n1705), .B1(n933), .Y(n3621) );
  OAI22XL U2457 ( .A0(n1680), .A1(n4068), .B0(n4063), .B1(n549), .Y(n3237) );
  OAI22XL U2458 ( .A0(n1679), .A1(n4023), .B0(n4018), .B1(n932), .Y(n3620) );
  OAI22XL U2459 ( .A0(n1679), .A1(n4067), .B0(n4063), .B1(n548), .Y(n3236) );
  OAI22XL U2460 ( .A0(n1678), .A1(n4023), .B0(n4018), .B1(n931), .Y(n3619) );
  OAI22XL U2461 ( .A0(n1678), .A1(n4064), .B0(n4063), .B1(n547), .Y(n3235) );
  OAI22XL U2462 ( .A0(n1677), .A1(n4023), .B0(n4018), .B1(n930), .Y(n3618) );
  OAI22XL U2463 ( .A0(n1677), .A1(n4065), .B0(n4063), .B1(n546), .Y(n3234) );
  OAI22XL U2464 ( .A0(n1676), .A1(n4023), .B0(n4018), .B1(n929), .Y(n3617) );
  OAI22XL U2465 ( .A0(n1676), .A1(n4068), .B0(n1698), .B1(n545), .Y(n3233) );
  OAI22XL U2466 ( .A0(n1675), .A1(n4023), .B0(n4018), .B1(n928), .Y(n3616) );
  OAI22XL U2467 ( .A0(n1675), .A1(n4067), .B0(n1698), .B1(n544), .Y(n3232) );
  OAI22XL U2468 ( .A0(n1674), .A1(n4023), .B0(n4018), .B1(n927), .Y(n3615) );
  OAI22XL U2469 ( .A0(n1674), .A1(n4065), .B0(n1698), .B1(n543), .Y(n3231) );
  OAI22XL U2470 ( .A0(n1673), .A1(n4023), .B0(n4018), .B1(n926), .Y(n3614) );
  OAI22XL U2471 ( .A0(n1673), .A1(n4066), .B0(n1698), .B1(n542), .Y(n3230) );
  OAI22XL U2472 ( .A0(n1618), .A1(n4023), .B0(n4020), .B1(n871), .Y(n3559) );
  OAI22XL U2473 ( .A0(n1618), .A1(n4072), .B0(n1338), .B1(n359), .Y(n3047) );
  OAI22XL U2474 ( .A0(n1617), .A1(n4022), .B0(n4021), .B1(n870), .Y(n3558) );
  OAI22XL U2475 ( .A0(n1617), .A1(n4072), .B0(n1339), .B1(n358), .Y(n3046) );
  OAI22XL U2476 ( .A0(n1616), .A1(n4024), .B0(n4017), .B1(n869), .Y(n3557) );
  OAI22XL U2477 ( .A0(n1616), .A1(n4072), .B0(n1338), .B1(n357), .Y(n3045) );
  OAI22XL U2478 ( .A0(n1615), .A1(n4023), .B0(n4017), .B1(n868), .Y(n3556) );
  OAI22XL U2479 ( .A0(n1615), .A1(n4073), .B0(n1339), .B1(n356), .Y(n3044) );
  OAI22XL U2480 ( .A0(n1614), .A1(n4022), .B0(n4017), .B1(n867), .Y(n3555) );
  OAI22XL U2481 ( .A0(n1614), .A1(n4077), .B0(n1338), .B1(n355), .Y(n3043) );
  OAI22XL U2482 ( .A0(n1613), .A1(n4024), .B0(n4017), .B1(n866), .Y(n3554) );
  OAI22XL U2483 ( .A0(n1613), .A1(n4072), .B0(n1339), .B1(n354), .Y(n3042) );
  OAI22XL U2484 ( .A0(n1612), .A1(n4023), .B0(n4017), .B1(n865), .Y(n3553) );
  OAI22XL U2485 ( .A0(n1612), .A1(n4072), .B0(n1338), .B1(n353), .Y(n3041) );
  OAI22XL U2486 ( .A0(n1545), .A1(n4023), .B0(n1705), .B1(n960), .Y(n3648) );
  OAI22XL U2487 ( .A0(n1545), .A1(n4075), .B0(n1338), .B1(n448), .Y(n3136) );
  OAI22XL U2488 ( .A0(n1544), .A1(n4022), .B0(n1705), .B1(n959), .Y(n3647) );
  OAI22XL U2489 ( .A0(n1544), .A1(n4074), .B0(n1339), .B1(n447), .Y(n3135) );
  OAI22XL U2490 ( .A0(n1543), .A1(n4024), .B0(n1705), .B1(n958), .Y(n3646) );
  OAI22XL U2491 ( .A0(n1543), .A1(n4073), .B0(n1338), .B1(n446), .Y(n3134) );
  OAI22XL U2492 ( .A0(n1542), .A1(n4028), .B0(n1705), .B1(n957), .Y(n3645) );
  OAI22XL U2493 ( .A0(n1542), .A1(n4077), .B0(n1339), .B1(n445), .Y(n3133) );
  OAI22XL U2494 ( .A0(n1541), .A1(n4028), .B0(n4017), .B1(n956), .Y(n3644) );
  OAI22XL U2495 ( .A0(n1541), .A1(n4072), .B0(n1338), .B1(n444), .Y(n3132) );
  OAI22XL U2496 ( .A0(n1540), .A1(n4023), .B0(n4017), .B1(n955), .Y(n3643) );
  OAI22XL U2497 ( .A0(n1540), .A1(n4075), .B0(n1339), .B1(n443), .Y(n3131) );
  OAI22XL U2498 ( .A0(n1602), .A1(n4028), .B0(n4021), .B1(n855), .Y(n3543) );
  OAI22XL U2499 ( .A0(n1601), .A1(n4028), .B0(n4016), .B1(n854), .Y(n3542) );
  OAI22XL U2500 ( .A0(n1600), .A1(n4028), .B0(n4016), .B1(n853), .Y(n3541) );
  OAI22XL U2501 ( .A0(n1599), .A1(n4022), .B0(n4016), .B1(n852), .Y(n3540) );
  OAI22XL U2502 ( .A0(n1598), .A1(n4028), .B0(n4016), .B1(n851), .Y(n3539) );
  OAI22XL U2503 ( .A0(n1597), .A1(n4023), .B0(n4016), .B1(n850), .Y(n3538) );
  OAI22XL U2504 ( .A0(n1596), .A1(n4022), .B0(n4016), .B1(n849), .Y(n3537) );
  OAI22XL U2505 ( .A0(n1595), .A1(n4024), .B0(n4016), .B1(n848), .Y(n3536) );
  OAI22XL U2506 ( .A0(n1594), .A1(n4026), .B0(n4016), .B1(n847), .Y(n3535) );
  OAI22XL U2507 ( .A0(n1593), .A1(n4026), .B0(n1706), .B1(n846), .Y(n3534) );
  OAI22XL U2508 ( .A0(n1592), .A1(n4025), .B0(n1706), .B1(n845), .Y(n3533) );
  OAI22XL U2509 ( .A0(n1591), .A1(n4027), .B0(n1706), .B1(n844), .Y(n3532) );
  OAI22XL U2510 ( .A0(n1590), .A1(n6), .B0(n1706), .B1(n843), .Y(n3531) );
  OAI22XL U2511 ( .A0(n1689), .A1(n4022), .B0(n1706), .B1(n942), .Y(n3630) );
  OAI22XL U2512 ( .A0(n1672), .A1(n4023), .B0(n4018), .B1(n925), .Y(n3613) );
  OAI22XL U2513 ( .A0(n1671), .A1(n4024), .B0(n4018), .B1(n924), .Y(n3612) );
  OAI22XL U2514 ( .A0(n1670), .A1(n4024), .B0(n4018), .B1(n923), .Y(n3611) );
  OAI22XL U2515 ( .A0(n1669), .A1(n4024), .B0(n4018), .B1(n922), .Y(n3610) );
  OAI22XL U2516 ( .A0(n1668), .A1(n4024), .B0(n4018), .B1(n921), .Y(n3609) );
  OAI22XL U2517 ( .A0(n1667), .A1(n4024), .B0(n4019), .B1(n920), .Y(n3608) );
  OAI22XL U2518 ( .A0(n1666), .A1(n4024), .B0(n4019), .B1(n919), .Y(n3607) );
  OAI22XL U2519 ( .A0(n1665), .A1(n4024), .B0(n4019), .B1(n918), .Y(n3606) );
  OAI22XL U2520 ( .A0(n1664), .A1(n4024), .B0(n4019), .B1(n917), .Y(n3605) );
  OAI22XL U2521 ( .A0(n1663), .A1(n4024), .B0(n4019), .B1(n916), .Y(n3604) );
  OAI22XL U2522 ( .A0(n1662), .A1(n4024), .B0(n4019), .B1(n915), .Y(n3603) );
  OAI22XL U2523 ( .A0(n1661), .A1(n4024), .B0(n4019), .B1(n914), .Y(n3602) );
  OAI22XL U2524 ( .A0(n1660), .A1(n4024), .B0(n4019), .B1(n913), .Y(n3601) );
  OAI22XL U2525 ( .A0(n1659), .A1(n4025), .B0(n4019), .B1(n912), .Y(n3600) );
  OAI22XL U2526 ( .A0(n1658), .A1(n4025), .B0(n4019), .B1(n911), .Y(n3599) );
  OAI22XL U2527 ( .A0(n1657), .A1(n4025), .B0(n4019), .B1(n910), .Y(n3598) );
  OAI22XL U2528 ( .A0(n1656), .A1(n4025), .B0(n4019), .B1(n909), .Y(n3597) );
  OAI22XL U2529 ( .A0(n1655), .A1(n4025), .B0(n4020), .B1(n908), .Y(n3596) );
  OAI22XL U2530 ( .A0(n1654), .A1(n4025), .B0(n4020), .B1(n907), .Y(n3595) );
  OAI22XL U2531 ( .A0(n1653), .A1(n4025), .B0(n4020), .B1(n906), .Y(n3594) );
  OAI22XL U2532 ( .A0(n1652), .A1(n4025), .B0(n4020), .B1(n905), .Y(n3593) );
  OAI22XL U2533 ( .A0(n1651), .A1(n4025), .B0(n4020), .B1(n904), .Y(n3592) );
  OAI22XL U2534 ( .A0(n1650), .A1(n4025), .B0(n4020), .B1(n903), .Y(n3591) );
  OAI22XL U2535 ( .A0(n1649), .A1(n4025), .B0(n4020), .B1(n902), .Y(n3590) );
  OAI22XL U2536 ( .A0(n1648), .A1(n4025), .B0(n4020), .B1(n901), .Y(n3589) );
  OAI22XL U2537 ( .A0(n1647), .A1(n4026), .B0(n4020), .B1(n900), .Y(n3588) );
  OAI22XL U2538 ( .A0(n1646), .A1(n4026), .B0(n4020), .B1(n899), .Y(n3587) );
  OAI22XL U2539 ( .A0(n1645), .A1(n4026), .B0(n4020), .B1(n898), .Y(n3586) );
  OAI22XL U2540 ( .A0(n1644), .A1(n4026), .B0(n4020), .B1(n897), .Y(n3585) );
  OAI22XL U2541 ( .A0(n1643), .A1(n4026), .B0(n4021), .B1(n896), .Y(n3584) );
  OAI22XL U2542 ( .A0(n1642), .A1(n4026), .B0(n4017), .B1(n895), .Y(n3583) );
  OAI22XL U2543 ( .A0(n1641), .A1(n4026), .B0(n4018), .B1(n894), .Y(n3582) );
  OAI22XL U2544 ( .A0(n1640), .A1(n4026), .B0(n4019), .B1(n893), .Y(n3581) );
  OAI22XL U2545 ( .A0(n1639), .A1(n4026), .B0(n4020), .B1(n892), .Y(n3580) );
  OAI22XL U2546 ( .A0(n1638), .A1(n4026), .B0(n4021), .B1(n891), .Y(n3579) );
  OAI22XL U2547 ( .A0(n1637), .A1(n4026), .B0(n4018), .B1(n890), .Y(n3578) );
  OAI22XL U2548 ( .A0(n1636), .A1(n4026), .B0(n4019), .B1(n889), .Y(n3577) );
  OAI22XL U2549 ( .A0(n1635), .A1(n4027), .B0(n4020), .B1(n888), .Y(n3576) );
  OAI22XL U2550 ( .A0(n1634), .A1(n4027), .B0(n4021), .B1(n887), .Y(n3575) );
  OAI22XL U2551 ( .A0(n1633), .A1(n4027), .B0(n4018), .B1(n886), .Y(n3574) );
  OAI22XL U2552 ( .A0(n1632), .A1(n4027), .B0(n4019), .B1(n885), .Y(n3573) );
  OAI22XL U2553 ( .A0(n1631), .A1(n4027), .B0(n4018), .B1(n884), .Y(n3572) );
  OAI22XL U2554 ( .A0(n1630), .A1(n4027), .B0(n4019), .B1(n883), .Y(n3571) );
  OAI22XL U2555 ( .A0(n1629), .A1(n4027), .B0(n4018), .B1(n882), .Y(n3570) );
  OAI22XL U2556 ( .A0(n1628), .A1(n4027), .B0(n4021), .B1(n881), .Y(n3569) );
  OAI22XL U2557 ( .A0(n1627), .A1(n4027), .B0(n4017), .B1(n880), .Y(n3568) );
  OAI22XL U2558 ( .A0(n1626), .A1(n4027), .B0(n4017), .B1(n879), .Y(n3567) );
  OAI22XL U2559 ( .A0(n1625), .A1(n4027), .B0(n4017), .B1(n878), .Y(n3566) );
  OAI22XL U2560 ( .A0(n1624), .A1(n4027), .B0(n4018), .B1(n877), .Y(n3565) );
  OAI22XL U2561 ( .A0(n1623), .A1(n4028), .B0(n4019), .B1(n876), .Y(n3564) );
  OAI22XL U2562 ( .A0(n1622), .A1(n4024), .B0(n4019), .B1(n875), .Y(n3563) );
  OAI22XL U2563 ( .A0(n1621), .A1(n4028), .B0(n4020), .B1(n874), .Y(n3562) );
  OAI22XL U2564 ( .A0(n1620), .A1(n4024), .B0(n4021), .B1(n873), .Y(n3561) );
  OAI22XL U2565 ( .A0(n1619), .A1(n4022), .B0(n4017), .B1(n872), .Y(n3560) );
  OAI22XL U2566 ( .A0(n1539), .A1(n4022), .B0(n4017), .B1(n954), .Y(n3642) );
  OAI22XL U2567 ( .A0(n1538), .A1(n4028), .B0(n1706), .B1(n953), .Y(n3641) );
  OAI22XL U2568 ( .A0(n1537), .A1(n4023), .B0(n1706), .B1(n952), .Y(n3640) );
  OAI22XL U2569 ( .A0(n1536), .A1(n4022), .B0(n1706), .B1(n951), .Y(n3639) );
  OAI22XL U2570 ( .A0(n1535), .A1(n4024), .B0(n1706), .B1(n950), .Y(n3638) );
  OAI22XL U2571 ( .A0(n1534), .A1(n4028), .B0(n1706), .B1(n949), .Y(n3637) );
  OAI22XL U2572 ( .A0(n1533), .A1(n4022), .B0(n1706), .B1(n948), .Y(n3636) );
  OAI22XL U2573 ( .A0(n1532), .A1(n4022), .B0(n4016), .B1(n947), .Y(n3635) );
  OAI22XL U2574 ( .A0(n1531), .A1(n4022), .B0(n4016), .B1(n946), .Y(n3634) );
  OAI22XL U2575 ( .A0(n1530), .A1(n4022), .B0(n4016), .B1(n945), .Y(n3633) );
  OAI22XL U2576 ( .A0(n1529), .A1(n4022), .B0(n4016), .B1(n944), .Y(n3632) );
  OAI22XL U2577 ( .A0(n1527), .A1(n4022), .B0(n4016), .B1(n943), .Y(n3631) );
  OAI221XL U2578 ( .A0(n1521), .A1(n4203), .B0(n1522), .B1(n4200), .C0(n1523), 
        .Y(proc_rdata[0]) );
  OA22X1 U2579 ( .A0(n1524), .A1(n4196), .B0(n1525), .B1(n4191), .Y(n1523) );
  OAI221XL U2580 ( .A0(n1466), .A1(n4202), .B0(n1467), .B1(n4199), .C0(n1468), 
        .Y(proc_rdata[1]) );
  OA22X1 U2581 ( .A0(n1469), .A1(n4194), .B0(n1470), .B1(n4192), .Y(n1468) );
  OAI221XL U2582 ( .A0(n1411), .A1(n4204), .B0(n1412), .B1(n4199), .C0(n1413), 
        .Y(proc_rdata[2]) );
  OA22X1 U2583 ( .A0(n1414), .A1(n4194), .B0(n1415), .B1(n4193), .Y(n1413) );
  OAI221XL U2584 ( .A0(n1396), .A1(n4204), .B0(n1397), .B1(n4198), .C0(n1398), 
        .Y(proc_rdata[3]) );
  OA22X1 U2585 ( .A0(n1399), .A1(n1368), .B0(n1400), .B1(n4193), .Y(n1398) );
  OAI221XL U2586 ( .A0(n1391), .A1(n4204), .B0(n1392), .B1(n4198), .C0(n1393), 
        .Y(proc_rdata[4]) );
  OA22X1 U2587 ( .A0(n1394), .A1(n1368), .B0(n1395), .B1(n4193), .Y(n1393) );
  OAI221XL U2588 ( .A0(n1386), .A1(n4204), .B0(n1387), .B1(n4198), .C0(n1388), 
        .Y(proc_rdata[5]) );
  OA22X1 U2589 ( .A0(n1389), .A1(n4196), .B0(n1390), .B1(n4192), .Y(n1388) );
  OAI221XL U2590 ( .A0(n1381), .A1(n4204), .B0(n1382), .B1(n4198), .C0(n1383), 
        .Y(proc_rdata[6]) );
  OA22X1 U2591 ( .A0(n1384), .A1(n1368), .B0(n1385), .B1(n4193), .Y(n1383) );
  OAI221XL U2592 ( .A0(n1376), .A1(n4204), .B0(n1377), .B1(n4198), .C0(n1378), 
        .Y(proc_rdata[7]) );
  OA22X1 U2593 ( .A0(n1379), .A1(n1368), .B0(n1380), .B1(n4193), .Y(n1378) );
  OAI221XL U2594 ( .A0(n1371), .A1(n4204), .B0(n1372), .B1(n4198), .C0(n1373), 
        .Y(proc_rdata[8]) );
  OA22X1 U2595 ( .A0(n1374), .A1(n1368), .B0(n1375), .B1(n4193), .Y(n1373) );
  OAI221XL U2596 ( .A0(n1362), .A1(n4203), .B0(n1364), .B1(n4199), .C0(n1366), 
        .Y(proc_rdata[9]) );
  OA22X1 U2597 ( .A0(n1367), .A1(n4196), .B0(n1369), .B1(n4192), .Y(n1366) );
  OAI221XL U2598 ( .A0(n1516), .A1(n4203), .B0(n1517), .B1(n4200), .C0(n1518), 
        .Y(proc_rdata[10]) );
  OA22X1 U2599 ( .A0(n1519), .A1(n4196), .B0(n1520), .B1(n4191), .Y(n1518) );
  OAI221XL U2600 ( .A0(n1511), .A1(n4203), .B0(n1512), .B1(n4200), .C0(n1513), 
        .Y(proc_rdata[11]) );
  OA22X1 U2601 ( .A0(n1514), .A1(n4196), .B0(n1515), .B1(n4191), .Y(n1513) );
  OAI221XL U2602 ( .A0(n1506), .A1(n4203), .B0(n1507), .B1(n4200), .C0(n1508), 
        .Y(proc_rdata[12]) );
  OA22X1 U2603 ( .A0(n1509), .A1(n4196), .B0(n1510), .B1(n4191), .Y(n1508) );
  OAI221XL U2604 ( .A0(n1501), .A1(n4201), .B0(n1502), .B1(n4200), .C0(n1503), 
        .Y(proc_rdata[13]) );
  OA22X1 U2605 ( .A0(n1504), .A1(n4196), .B0(n1505), .B1(n4191), .Y(n1503) );
  OAI221XL U2606 ( .A0(n1496), .A1(n4201), .B0(n1497), .B1(n4200), .C0(n1498), 
        .Y(proc_rdata[14]) );
  OA22X1 U2607 ( .A0(n1499), .A1(n4196), .B0(n1500), .B1(n4191), .Y(n1498) );
  OAI221XL U2608 ( .A0(n1491), .A1(n9), .B0(n1492), .B1(n4200), .C0(n1493), 
        .Y(proc_rdata[15]) );
  OA22X1 U2609 ( .A0(n1494), .A1(n4195), .B0(n1495), .B1(n4193), .Y(n1493) );
  OAI221XL U2610 ( .A0(n1486), .A1(n4203), .B0(n1487), .B1(n4200), .C0(n1488), 
        .Y(proc_rdata[16]) );
  OA22X1 U2611 ( .A0(n1489), .A1(n4194), .B0(n1490), .B1(n4191), .Y(n1488) );
  OAI221XL U2612 ( .A0(n1481), .A1(n4201), .B0(n1482), .B1(n4200), .C0(n1483), 
        .Y(proc_rdata[17]) );
  OA22X1 U2613 ( .A0(n1484), .A1(n4195), .B0(n1485), .B1(n4191), .Y(n1483) );
  OAI221XL U2614 ( .A0(n1476), .A1(n4201), .B0(n1477), .B1(n4200), .C0(n1478), 
        .Y(proc_rdata[18]) );
  OA22X1 U2615 ( .A0(n1479), .A1(n4196), .B0(n1480), .B1(n4191), .Y(n1478) );
  OAI221XL U2616 ( .A0(n1471), .A1(n4201), .B0(n1472), .B1(n4199), .C0(n1473), 
        .Y(proc_rdata[19]) );
  OA22X1 U2617 ( .A0(n1474), .A1(n4194), .B0(n1475), .B1(n16), .Y(n1473) );
  OAI221XL U2618 ( .A0(n1461), .A1(n9), .B0(n1462), .B1(n4199), .C0(n1463), 
        .Y(proc_rdata[20]) );
  OA22X1 U2619 ( .A0(n1464), .A1(n4196), .B0(n1465), .B1(n16), .Y(n1463) );
  OAI221XL U2620 ( .A0(n1456), .A1(n9), .B0(n1457), .B1(n4199), .C0(n1458), 
        .Y(proc_rdata[21]) );
  OA22X1 U2621 ( .A0(n1459), .A1(n4194), .B0(n1460), .B1(n16), .Y(n1458) );
  OAI221XL U2622 ( .A0(n1451), .A1(n4203), .B0(n1452), .B1(n4199), .C0(n1453), 
        .Y(proc_rdata[22]) );
  OA22X1 U2623 ( .A0(n1454), .A1(n4194), .B0(n1455), .B1(n4192), .Y(n1453) );
  OAI221XL U2624 ( .A0(n1446), .A1(n4202), .B0(n1447), .B1(n4199), .C0(n1448), 
        .Y(proc_rdata[23]) );
  OA22X1 U2625 ( .A0(n1449), .A1(n4195), .B0(n1450), .B1(n4192), .Y(n1448) );
  OAI221XL U2626 ( .A0(n1441), .A1(n9), .B0(n1442), .B1(n4199), .C0(n1443), 
        .Y(proc_rdata[24]) );
  OA22X1 U2627 ( .A0(n1444), .A1(n4196), .B0(n1445), .B1(n16), .Y(n1443) );
  OAI221XL U2628 ( .A0(n1436), .A1(n4204), .B0(n1437), .B1(n4199), .C0(n1438), 
        .Y(proc_rdata[25]) );
  OA22X1 U2629 ( .A0(n1439), .A1(n4195), .B0(n1440), .B1(n4193), .Y(n1438) );
  OAI221XL U2630 ( .A0(n1431), .A1(n9), .B0(n1432), .B1(n4199), .C0(n1433), 
        .Y(proc_rdata[26]) );
  OA22X1 U2631 ( .A0(n1434), .A1(n4194), .B0(n1435), .B1(n16), .Y(n1433) );
  OAI221XL U2632 ( .A0(n1426), .A1(n4202), .B0(n1427), .B1(n4199), .C0(n1428), 
        .Y(proc_rdata[27]) );
  OA22X1 U2633 ( .A0(n1429), .A1(n4195), .B0(n1430), .B1(n4192), .Y(n1428) );
  OAI221XL U2634 ( .A0(n1421), .A1(n4204), .B0(n1422), .B1(n4199), .C0(n1423), 
        .Y(proc_rdata[28]) );
  OA22X1 U2635 ( .A0(n1424), .A1(n4195), .B0(n1425), .B1(n16), .Y(n1423) );
  OAI221XL U2636 ( .A0(n1416), .A1(n4204), .B0(n1417), .B1(n4199), .C0(n1418), 
        .Y(proc_rdata[29]) );
  OA22X1 U2637 ( .A0(n1419), .A1(n4195), .B0(n1420), .B1(n4193), .Y(n1418) );
  OAI221XL U2638 ( .A0(n1406), .A1(n9), .B0(n1407), .B1(n4199), .C0(n1408), 
        .Y(proc_rdata[30]) );
  OA22X1 U2639 ( .A0(n1409), .A1(n4195), .B0(n1410), .B1(n4191), .Y(n1408) );
  OAI221XL U2640 ( .A0(n1401), .A1(n4204), .B0(n1402), .B1(n4199), .C0(n1403), 
        .Y(proc_rdata[31]) );
  OA22X1 U2641 ( .A0(n1404), .A1(n4195), .B0(n1405), .B1(n4193), .Y(n1403) );
  NAND2XL U2642 ( .A(proc_write), .B(n4353), .Y(n1576) );
  INVXL U2643 ( .A(proc_addr_0), .Y(n4354) );
  INVXL U2644 ( .A(proc_addr_1), .Y(n4355) );
  OAI22XL U2645 ( .A0(n64), .A1(n1565), .B0(n4349), .B1(n1566), .Y(n3992) );
  AOI2BB1XL U2646 ( .A0N(n1360), .A1N(n4351), .B0(n4419), .Y(n1566) );
  CLKINVX1 U2647 ( .A(n1567), .Y(n4351) );
  OAI22XL U2648 ( .A0(n4131), .A1(n288), .B0(n4144), .B1(n160), .Y(n2413) );
  OAI22XL U2649 ( .A0(n4116), .A1(n544), .B0(n4125), .B1(n416), .Y(n2414) );
  OAI22XL U2650 ( .A0(n1696), .A1(n800), .B0(n1370), .B1(n672), .Y(n2411) );
  OAI22XL U2651 ( .A0(n4135), .A1(n287), .B0(n4144), .B1(n159), .Y(n2409) );
  OAI22XL U2652 ( .A0(n4116), .A1(n543), .B0(n4127), .B1(n415), .Y(n2410) );
  OAI22XL U2653 ( .A0(n1696), .A1(n799), .B0(n1370), .B1(n671), .Y(n2407) );
  OAI22XL U2654 ( .A0(n4137), .A1(n286), .B0(n4144), .B1(n158), .Y(n2405) );
  OAI22XL U2655 ( .A0(n4116), .A1(n542), .B0(n4125), .B1(n414), .Y(n2406) );
  OAI22XL U2656 ( .A0(n1696), .A1(n798), .B0(n1370), .B1(n670), .Y(n2403) );
  OAI22XL U2657 ( .A0(n4133), .A1(n285), .B0(n4144), .B1(n157), .Y(n2401) );
  OAI22XL U2658 ( .A0(n4116), .A1(n541), .B0(n4123), .B1(n413), .Y(n2402) );
  OAI22XL U2659 ( .A0(n1696), .A1(n797), .B0(n1370), .B1(n669), .Y(n2399) );
  OAI22XL U2660 ( .A0(n4133), .A1(n284), .B0(n4144), .B1(n156), .Y(n2397) );
  OAI22XL U2661 ( .A0(n4116), .A1(n540), .B0(n4123), .B1(n412), .Y(n2398) );
  OAI22XL U2662 ( .A0(n1696), .A1(n796), .B0(n1370), .B1(n668), .Y(n2395) );
  OAI22XL U2663 ( .A0(n4133), .A1(n283), .B0(n4144), .B1(n155), .Y(n2393) );
  OAI22XL U2664 ( .A0(n4116), .A1(n539), .B0(n4123), .B1(n411), .Y(n2394) );
  OAI22XL U2665 ( .A0(n1696), .A1(n795), .B0(n1370), .B1(n667), .Y(n2391) );
  OAI22XL U2666 ( .A0(n4135), .A1(n282), .B0(n4144), .B1(n154), .Y(n2389) );
  OAI22XL U2667 ( .A0(n4116), .A1(n538), .B0(n4127), .B1(n410), .Y(n2390) );
  OAI22XL U2668 ( .A0(n1696), .A1(n794), .B0(n1370), .B1(n666), .Y(n2387) );
  OAI22XL U2669 ( .A0(n4137), .A1(n281), .B0(n4144), .B1(n153), .Y(n2385) );
  OAI22XL U2670 ( .A0(n4116), .A1(n537), .B0(n4125), .B1(n409), .Y(n2386) );
  OAI22XL U2671 ( .A0(n1696), .A1(n793), .B0(n1370), .B1(n665), .Y(n2383) );
  OAI22XL U2672 ( .A0(n4136), .A1(n280), .B0(n4144), .B1(n152), .Y(n2377) );
  OAI22XL U2673 ( .A0(n4116), .A1(n536), .B0(n4126), .B1(n408), .Y(n2378) );
  OAI22XL U2674 ( .A0(n1696), .A1(n792), .B0(n1370), .B1(n664), .Y(n2375) );
  OAI22XL U2675 ( .A0(n4134), .A1(n279), .B0(n4144), .B1(n151), .Y(n2373) );
  OAI22XL U2676 ( .A0(n4116), .A1(n535), .B0(n4124), .B1(n407), .Y(n2374) );
  OAI22XL U2677 ( .A0(n1696), .A1(n791), .B0(n1370), .B1(n663), .Y(n2371) );
  OAI22XL U2678 ( .A0(n4135), .A1(n278), .B0(n4143), .B1(n150), .Y(n2369) );
  OAI22XL U2679 ( .A0(n4115), .A1(n534), .B0(n4125), .B1(n406), .Y(n2370) );
  OAI22XL U2680 ( .A0(n1695), .A1(n790), .B0(n1358), .B1(n662), .Y(n2367) );
  OAI22XL U2681 ( .A0(n4135), .A1(n277), .B0(n4143), .B1(n149), .Y(n2365) );
  OAI22XL U2682 ( .A0(n4115), .A1(n533), .B0(n4125), .B1(n405), .Y(n2366) );
  OAI22XL U2683 ( .A0(n1695), .A1(n789), .B0(n1370), .B1(n661), .Y(n2363) );
  OAI22XL U2684 ( .A0(n4135), .A1(n276), .B0(n4143), .B1(n148), .Y(n2361) );
  OAI22XL U2685 ( .A0(n4115), .A1(n532), .B0(n4125), .B1(n404), .Y(n2362) );
  OAI22XL U2686 ( .A0(n1695), .A1(n788), .B0(n1358), .B1(n660), .Y(n2359) );
  OAI22XL U2687 ( .A0(n4135), .A1(n275), .B0(n4143), .B1(n147), .Y(n2357) );
  OAI22XL U2688 ( .A0(n4115), .A1(n531), .B0(n4125), .B1(n403), .Y(n2358) );
  OAI22XL U2689 ( .A0(n1695), .A1(n787), .B0(n1358), .B1(n659), .Y(n2355) );
  OAI22XL U2690 ( .A0(n4135), .A1(n274), .B0(n4143), .B1(n146), .Y(n2353) );
  OAI22XL U2691 ( .A0(n4115), .A1(n530), .B0(n4125), .B1(n402), .Y(n2354) );
  OAI22XL U2692 ( .A0(n1695), .A1(n786), .B0(n1358), .B1(n658), .Y(n2351) );
  OAI22XL U2693 ( .A0(n4135), .A1(n273), .B0(n4143), .B1(n145), .Y(n2349) );
  OAI22XL U2694 ( .A0(n4115), .A1(n529), .B0(n4125), .B1(n401), .Y(n2350) );
  OAI22XL U2695 ( .A0(n1695), .A1(n785), .B0(n1358), .B1(n657), .Y(n2347) );
  OAI22XL U2696 ( .A0(n4135), .A1(n272), .B0(n4143), .B1(n144), .Y(n2345) );
  OAI22XL U2697 ( .A0(n4115), .A1(n528), .B0(n4125), .B1(n400), .Y(n2346) );
  OAI22XL U2698 ( .A0(n1695), .A1(n784), .B0(n1358), .B1(n656), .Y(n2343) );
  OAI22XL U2699 ( .A0(n4135), .A1(n271), .B0(n4143), .B1(n143), .Y(n2341) );
  OAI22XL U2700 ( .A0(n4115), .A1(n527), .B0(n4125), .B1(n399), .Y(n2342) );
  OAI22XL U2701 ( .A0(n1695), .A1(n783), .B0(n1359), .B1(n655), .Y(n2339) );
  OAI22XL U2702 ( .A0(n4135), .A1(n270), .B0(n4143), .B1(n142), .Y(n2333) );
  OAI22XL U2703 ( .A0(n4115), .A1(n526), .B0(n4125), .B1(n398), .Y(n2334) );
  OAI22XL U2704 ( .A0(n1695), .A1(n782), .B0(n1359), .B1(n654), .Y(n2331) );
  OAI22XL U2705 ( .A0(n4135), .A1(n269), .B0(n4143), .B1(n141), .Y(n2329) );
  OAI22XL U2706 ( .A0(n4115), .A1(n525), .B0(n4125), .B1(n397), .Y(n2330) );
  OAI22XL U2707 ( .A0(n1695), .A1(n781), .B0(n1359), .B1(n653), .Y(n2327) );
  OAI22XL U2708 ( .A0(n4135), .A1(n268), .B0(n4143), .B1(n140), .Y(n2325) );
  OAI22XL U2709 ( .A0(n4115), .A1(n524), .B0(n4125), .B1(n396), .Y(n2326) );
  OAI22XL U2710 ( .A0(n1695), .A1(n780), .B0(n1359), .B1(n652), .Y(n2323) );
  OAI22XL U2711 ( .A0(n4135), .A1(n267), .B0(n4143), .B1(n139), .Y(n2321) );
  OAI22XL U2712 ( .A0(n4115), .A1(n523), .B0(n4125), .B1(n395), .Y(n2322) );
  OAI22XL U2713 ( .A0(n1695), .A1(n779), .B0(n1359), .B1(n651), .Y(n2319) );
  OAI22XL U2714 ( .A0(n4135), .A1(n266), .B0(n4143), .B1(n138), .Y(n2317) );
  OAI22XL U2715 ( .A0(n4115), .A1(n522), .B0(n4125), .B1(n394), .Y(n2318) );
  OAI22XL U2716 ( .A0(n1695), .A1(n778), .B0(n1359), .B1(n650), .Y(n2315) );
  OAI22XL U2717 ( .A0(n4135), .A1(n265), .B0(n4143), .B1(n137), .Y(n2313) );
  OAI22XL U2718 ( .A0(n4115), .A1(n521), .B0(n4125), .B1(n393), .Y(n2314) );
  OAI22XL U2719 ( .A0(n1695), .A1(n777), .B0(n1363), .B1(n649), .Y(n2311) );
  OAI22XL U2720 ( .A0(n4135), .A1(n264), .B0(n4143), .B1(n136), .Y(n2309) );
  OAI22XL U2721 ( .A0(n4115), .A1(n520), .B0(n4125), .B1(n392), .Y(n2310) );
  OAI22XL U2722 ( .A0(n1695), .A1(n776), .B0(n1358), .B1(n648), .Y(n2307) );
  OAI22XL U2723 ( .A0(n4135), .A1(n263), .B0(n4143), .B1(n135), .Y(n2305) );
  OAI22XL U2724 ( .A0(n4115), .A1(n519), .B0(n4125), .B1(n391), .Y(n2306) );
  OAI22XL U2725 ( .A0(n1695), .A1(n775), .B0(n1358), .B1(n647), .Y(n2303) );
  OAI22XL U2726 ( .A0(n4134), .A1(n262), .B0(n4142), .B1(n134), .Y(n2301) );
  OAI22XL U2727 ( .A0(n4114), .A1(n518), .B0(n4124), .B1(n390), .Y(n2302) );
  OAI22XL U2728 ( .A0(n4359), .A1(n774), .B0(n1365), .B1(n646), .Y(n2299) );
  OAI22XL U2729 ( .A0(n4134), .A1(n261), .B0(n4142), .B1(n133), .Y(n2297) );
  OAI22XL U2730 ( .A0(n4114), .A1(n517), .B0(n4124), .B1(n389), .Y(n2298) );
  OAI22XL U2731 ( .A0(n1558), .A1(n773), .B0(n1365), .B1(n645), .Y(n2295) );
  OAI22XL U2732 ( .A0(n4134), .A1(n260), .B0(n4142), .B1(n132), .Y(n2289) );
  OAI22XL U2733 ( .A0(n4114), .A1(n516), .B0(n4124), .B1(n388), .Y(n2290) );
  OAI22XL U2734 ( .A0(n1558), .A1(n772), .B0(n1365), .B1(n644), .Y(n2287) );
  OAI22XL U2735 ( .A0(n4134), .A1(n259), .B0(n4142), .B1(n131), .Y(n2285) );
  OAI22XL U2736 ( .A0(n4114), .A1(n515), .B0(n4124), .B1(n387), .Y(n2286) );
  OAI22XL U2737 ( .A0(n1558), .A1(n771), .B0(n1365), .B1(n643), .Y(n2283) );
  OAI22XL U2738 ( .A0(n4134), .A1(n258), .B0(n4142), .B1(n130), .Y(n2281) );
  OAI22XL U2739 ( .A0(n4114), .A1(n514), .B0(n4124), .B1(n386), .Y(n2282) );
  OAI22XL U2740 ( .A0(n1558), .A1(n770), .B0(n1365), .B1(n642), .Y(n2279) );
  OAI22XL U2741 ( .A0(n4134), .A1(n257), .B0(n4142), .B1(n129), .Y(n2277) );
  OAI22XL U2742 ( .A0(n4114), .A1(n513), .B0(n4124), .B1(n385), .Y(n2278) );
  OAI22XL U2743 ( .A0(n1558), .A1(n769), .B0(n1365), .B1(n641), .Y(n2275) );
  OAI22XL U2744 ( .A0(n4134), .A1(n256), .B0(n4142), .B1(n128), .Y(n2273) );
  OAI22XL U2745 ( .A0(n4114), .A1(n512), .B0(n4124), .B1(n384), .Y(n2274) );
  OAI22XL U2746 ( .A0(n1696), .A1(n768), .B0(n1365), .B1(n640), .Y(n2271) );
  OAI22XL U2747 ( .A0(n4134), .A1(n255), .B0(n4142), .B1(n127), .Y(n2269) );
  OAI22XL U2748 ( .A0(n4114), .A1(n511), .B0(n4124), .B1(n383), .Y(n2270) );
  OAI22XL U2749 ( .A0(n1695), .A1(n767), .B0(n1365), .B1(n639), .Y(n2267) );
  OAI22XL U2750 ( .A0(n4134), .A1(n254), .B0(n4142), .B1(n126), .Y(n2265) );
  OAI22XL U2751 ( .A0(n4114), .A1(n510), .B0(n4124), .B1(n382), .Y(n2266) );
  OAI22XL U2752 ( .A0(n1697), .A1(n766), .B0(n1365), .B1(n638), .Y(n2263) );
  OAI22XL U2753 ( .A0(n4134), .A1(n253), .B0(n4142), .B1(n125), .Y(n2261) );
  OAI22XL U2754 ( .A0(n4114), .A1(n509), .B0(n4124), .B1(n381), .Y(n2262) );
  OAI22XL U2755 ( .A0(n1580), .A1(n765), .B0(n1365), .B1(n637), .Y(n2259) );
  OAI22XL U2756 ( .A0(n4134), .A1(n252), .B0(n4142), .B1(n124), .Y(n2257) );
  OAI22XL U2757 ( .A0(n4114), .A1(n508), .B0(n4124), .B1(n380), .Y(n2258) );
  OAI22XL U2758 ( .A0(n1558), .A1(n764), .B0(n1365), .B1(n636), .Y(n2255) );
  OAI22XL U2759 ( .A0(n4134), .A1(n251), .B0(n4142), .B1(n123), .Y(n2253) );
  OAI22XL U2760 ( .A0(n4114), .A1(n507), .B0(n4124), .B1(n379), .Y(n2254) );
  OAI22XL U2761 ( .A0(n1558), .A1(n763), .B0(n1365), .B1(n635), .Y(n2251) );
  OAI22XL U2762 ( .A0(n4134), .A1(n250), .B0(n4142), .B1(n122), .Y(n2245) );
  OAI22XL U2763 ( .A0(n4114), .A1(n506), .B0(n4124), .B1(n378), .Y(n2246) );
  OAI22XL U2764 ( .A0(n1558), .A1(n762), .B0(n1365), .B1(n634), .Y(n2243) );
  OAI22XL U2765 ( .A0(n4134), .A1(n249), .B0(n4142), .B1(n121), .Y(n2241) );
  OAI22XL U2766 ( .A0(n4114), .A1(n505), .B0(n4124), .B1(n377), .Y(n2242) );
  OAI22XL U2767 ( .A0(n4359), .A1(n761), .B0(n1365), .B1(n633), .Y(n2239) );
  OAI22XL U2768 ( .A0(n4134), .A1(n248), .B0(n4142), .B1(n120), .Y(n2237) );
  OAI22XL U2769 ( .A0(n4114), .A1(n504), .B0(n4124), .B1(n376), .Y(n2238) );
  OAI22XL U2770 ( .A0(n4359), .A1(n760), .B0(n1365), .B1(n632), .Y(n2235) );
  OAI22XL U2771 ( .A0(n4134), .A1(n247), .B0(n4142), .B1(n119), .Y(n2233) );
  OAI22XL U2772 ( .A0(n4114), .A1(n503), .B0(n4124), .B1(n375), .Y(n2234) );
  OAI22XL U2773 ( .A0(n4359), .A1(n759), .B0(n1365), .B1(n631), .Y(n2231) );
  OAI22XL U2774 ( .A0(n4133), .A1(n246), .B0(n4148), .B1(n118), .Y(n2229) );
  OAI22XL U2775 ( .A0(n4113), .A1(n502), .B0(n4123), .B1(n374), .Y(n2230) );
  OAI22XL U2776 ( .A0(n1693), .A1(n758), .B0(n4357), .B1(n630), .Y(n2227) );
  OAI22XL U2777 ( .A0(n4133), .A1(n245), .B0(n4147), .B1(n117), .Y(n2225) );
  OAI22XL U2778 ( .A0(n4113), .A1(n501), .B0(n4123), .B1(n373), .Y(n2226) );
  OAI22XL U2779 ( .A0(n1693), .A1(n757), .B0(n1359), .B1(n629), .Y(n2223) );
  OAI22XL U2780 ( .A0(n4133), .A1(n244), .B0(n4146), .B1(n116), .Y(n2221) );
  OAI22XL U2781 ( .A0(n4113), .A1(n500), .B0(n4123), .B1(n372), .Y(n2222) );
  OAI22XL U2782 ( .A0(n1693), .A1(n756), .B0(n1359), .B1(n628), .Y(n2219) );
  OAI22XL U2783 ( .A0(n4133), .A1(n243), .B0(n4145), .B1(n115), .Y(n2217) );
  OAI22XL U2784 ( .A0(n4113), .A1(n499), .B0(n4123), .B1(n371), .Y(n2218) );
  OAI22XL U2785 ( .A0(n1693), .A1(n755), .B0(n1359), .B1(n627), .Y(n2215) );
  OAI22XL U2786 ( .A0(n4133), .A1(n242), .B0(n4143), .B1(n114), .Y(n2213) );
  OAI22XL U2787 ( .A0(n4113), .A1(n498), .B0(n4123), .B1(n370), .Y(n2214) );
  OAI22XL U2788 ( .A0(n1693), .A1(n754), .B0(n1359), .B1(n626), .Y(n2211) );
  OAI22XL U2789 ( .A0(n4133), .A1(n241), .B0(n4144), .B1(n113), .Y(n2209) );
  OAI22XL U2790 ( .A0(n4113), .A1(n497), .B0(n4123), .B1(n369), .Y(n2210) );
  OAI22XL U2791 ( .A0(n1693), .A1(n753), .B0(n1359), .B1(n625), .Y(n2207) );
  OAI22XL U2792 ( .A0(n4133), .A1(n240), .B0(n4142), .B1(n112), .Y(n2201) );
  OAI22XL U2793 ( .A0(n4113), .A1(n496), .B0(n4123), .B1(n368), .Y(n2202) );
  OAI22XL U2794 ( .A0(n1693), .A1(n752), .B0(n1359), .B1(n624), .Y(n2199) );
  OAI22XL U2795 ( .A0(n4133), .A1(n239), .B0(n4146), .B1(n111), .Y(n2197) );
  OAI22XL U2796 ( .A0(n4113), .A1(n495), .B0(n4123), .B1(n367), .Y(n2198) );
  OAI22XL U2797 ( .A0(n1693), .A1(n751), .B0(n1359), .B1(n623), .Y(n2195) );
  OAI22XL U2798 ( .A0(n4133), .A1(n238), .B0(n4145), .B1(n110), .Y(n2193) );
  OAI22XL U2799 ( .A0(n4113), .A1(n494), .B0(n4123), .B1(n366), .Y(n2194) );
  OAI22XL U2800 ( .A0(n1693), .A1(n750), .B0(n1359), .B1(n622), .Y(n2191) );
  OAI22XL U2801 ( .A0(n4133), .A1(n237), .B0(n4143), .B1(n109), .Y(n2189) );
  OAI22XL U2802 ( .A0(n4113), .A1(n493), .B0(n4123), .B1(n365), .Y(n2190) );
  OAI22XL U2803 ( .A0(n1693), .A1(n749), .B0(n4357), .B1(n621), .Y(n2187) );
  OAI22XL U2804 ( .A0(n4133), .A1(n236), .B0(n4144), .B1(n108), .Y(n2185) );
  OAI22XL U2805 ( .A0(n4113), .A1(n492), .B0(n4123), .B1(n364), .Y(n2186) );
  OAI22XL U2806 ( .A0(n1693), .A1(n748), .B0(n1359), .B1(n620), .Y(n2183) );
  OAI22XL U2807 ( .A0(n4133), .A1(n235), .B0(n4142), .B1(n107), .Y(n2181) );
  OAI22XL U2808 ( .A0(n4113), .A1(n491), .B0(n4123), .B1(n363), .Y(n2182) );
  OAI22XL U2809 ( .A0(n1693), .A1(n747), .B0(n4357), .B1(n619), .Y(n2179) );
  OAI22XL U2810 ( .A0(n4133), .A1(n234), .B0(n4148), .B1(n106), .Y(n2177) );
  OAI22XL U2811 ( .A0(n4113), .A1(n490), .B0(n4123), .B1(n362), .Y(n2178) );
  OAI22XL U2812 ( .A0(n1693), .A1(n746), .B0(n4357), .B1(n618), .Y(n2175) );
  OAI22XL U2813 ( .A0(n4133), .A1(n233), .B0(n4147), .B1(n105), .Y(n2173) );
  OAI22XL U2814 ( .A0(n4113), .A1(n489), .B0(n4123), .B1(n361), .Y(n2174) );
  OAI22XL U2815 ( .A0(n1693), .A1(n745), .B0(n1359), .B1(n617), .Y(n2171) );
  OAI22XL U2816 ( .A0(n4133), .A1(n232), .B0(n4148), .B1(n104), .Y(n2169) );
  OAI22XL U2817 ( .A0(n4113), .A1(n488), .B0(n4123), .B1(n360), .Y(n2170) );
  OAI22XL U2818 ( .A0(n1693), .A1(n744), .B0(n1359), .B1(n616), .Y(n2167) );
  OAI22XL U2819 ( .A0(n4132), .A1(n231), .B0(n4141), .B1(n103), .Y(n2165) );
  OAI22XL U2820 ( .A0(n4112), .A1(n487), .B0(n4122), .B1(n359), .Y(n2166) );
  OAI22XL U2821 ( .A0(n1580), .A1(n743), .B0(n1363), .B1(n615), .Y(n2163) );
  OAI22XL U2822 ( .A0(n4132), .A1(n230), .B0(n4141), .B1(n102), .Y(n2157) );
  OAI22XL U2823 ( .A0(n4112), .A1(n486), .B0(n4122), .B1(n358), .Y(n2158) );
  OAI22XL U2824 ( .A0(n1580), .A1(n742), .B0(n1363), .B1(n614), .Y(n2155) );
  OAI22XL U2825 ( .A0(n4132), .A1(n229), .B0(n4141), .B1(n101), .Y(n2153) );
  OAI22XL U2826 ( .A0(n4112), .A1(n485), .B0(n4122), .B1(n357), .Y(n2154) );
  OAI22XL U2827 ( .A0(n1580), .A1(n741), .B0(n1363), .B1(n613), .Y(n2151) );
  OAI22XL U2828 ( .A0(n4132), .A1(n228), .B0(n4141), .B1(n100), .Y(n2149) );
  OAI22XL U2829 ( .A0(n4112), .A1(n484), .B0(n4122), .B1(n356), .Y(n2150) );
  OAI22XL U2830 ( .A0(n1580), .A1(n740), .B0(n1363), .B1(n612), .Y(n2147) );
  OAI22XL U2831 ( .A0(n4132), .A1(n227), .B0(n4141), .B1(n99), .Y(n2145) );
  OAI22XL U2832 ( .A0(n4112), .A1(n483), .B0(n4122), .B1(n355), .Y(n2146) );
  OAI22XL U2833 ( .A0(n1580), .A1(n739), .B0(n1363), .B1(n611), .Y(n2143) );
  OAI22XL U2834 ( .A0(n4132), .A1(n226), .B0(n4141), .B1(n98), .Y(n2141) );
  OAI22XL U2835 ( .A0(n4112), .A1(n482), .B0(n4122), .B1(n354), .Y(n2142) );
  OAI22XL U2836 ( .A0(n1580), .A1(n738), .B0(n1363), .B1(n610), .Y(n2139) );
  OAI22XL U2837 ( .A0(n4132), .A1(n225), .B0(n4141), .B1(n97), .Y(n2137) );
  OAI22XL U2838 ( .A0(n4112), .A1(n481), .B0(n4122), .B1(n353), .Y(n2138) );
  OAI22XL U2839 ( .A0(n1580), .A1(n737), .B0(n1363), .B1(n609), .Y(n2135) );
  OAI22XL U2840 ( .A0(n4132), .A1(n224), .B0(n4141), .B1(n96), .Y(n2133) );
  OAI22XL U2841 ( .A0(n4112), .A1(n480), .B0(n4122), .B1(n352), .Y(n2134) );
  OAI22XL U2842 ( .A0(n1580), .A1(n736), .B0(n1363), .B1(n608), .Y(n2131) );
  OAI22XL U2843 ( .A0(n4132), .A1(n223), .B0(n4141), .B1(n95), .Y(n2129) );
  OAI22XL U2844 ( .A0(n4112), .A1(n479), .B0(n4122), .B1(n351), .Y(n2130) );
  OAI22XL U2845 ( .A0(n1580), .A1(n735), .B0(n1363), .B1(n607), .Y(n2127) );
  OAI22XL U2846 ( .A0(n4132), .A1(n222), .B0(n4141), .B1(n94), .Y(n2125) );
  OAI22XL U2847 ( .A0(n4112), .A1(n478), .B0(n4122), .B1(n350), .Y(n2126) );
  OAI22XL U2848 ( .A0(n1580), .A1(n734), .B0(n1363), .B1(n606), .Y(n2123) );
  OAI22XL U2849 ( .A0(n4132), .A1(n221), .B0(n4141), .B1(n93), .Y(n2121) );
  OAI22XL U2850 ( .A0(n4112), .A1(n477), .B0(n4122), .B1(n349), .Y(n2122) );
  OAI22XL U2851 ( .A0(n1580), .A1(n733), .B0(n1363), .B1(n605), .Y(n2119) );
  OAI22XL U2852 ( .A0(n4137), .A1(n220), .B0(n4147), .B1(n92), .Y(n2621) );
  OAI22XL U2853 ( .A0(n4118), .A1(n476), .B0(n4127), .B1(n348), .Y(n2622) );
  OAI22XL U2854 ( .A0(n1701), .A1(n732), .B0(n1546), .B1(n604), .Y(n2619) );
  OAI22XL U2855 ( .A0(n4137), .A1(n219), .B0(n4147), .B1(n91), .Y(n2617) );
  OAI22XL U2856 ( .A0(n4118), .A1(n475), .B0(n4127), .B1(n347), .Y(n2618) );
  OAI22XL U2857 ( .A0(n1701), .A1(n731), .B0(n1546), .B1(n603), .Y(n2615) );
  OAI22XL U2858 ( .A0(n4137), .A1(n218), .B0(n4147), .B1(n90), .Y(n2613) );
  OAI22XL U2859 ( .A0(n4118), .A1(n474), .B0(n4127), .B1(n346), .Y(n2614) );
  OAI22XL U2860 ( .A0(n1701), .A1(n730), .B0(n1546), .B1(n602), .Y(n2611) );
  OAI22XL U2861 ( .A0(n4137), .A1(n217), .B0(n4147), .B1(n89), .Y(n2609) );
  OAI22XL U2862 ( .A0(n4118), .A1(n473), .B0(n4127), .B1(n345), .Y(n2610) );
  OAI22XL U2863 ( .A0(n1701), .A1(n729), .B0(n1546), .B1(n601), .Y(n2607) );
  OAI22XL U2864 ( .A0(n4137), .A1(n216), .B0(n4147), .B1(n88), .Y(n2605) );
  OAI22XL U2865 ( .A0(n4118), .A1(n472), .B0(n4127), .B1(n344), .Y(n2606) );
  OAI22XL U2866 ( .A0(n1701), .A1(n728), .B0(n1546), .B1(n600), .Y(n2603) );
  OAI22XL U2867 ( .A0(n4137), .A1(n215), .B0(n4147), .B1(n87), .Y(n2601) );
  OAI22XL U2868 ( .A0(n4118), .A1(n471), .B0(n4127), .B1(n343), .Y(n2602) );
  OAI22XL U2869 ( .A0(n1701), .A1(n727), .B0(n1546), .B1(n599), .Y(n2599) );
  OAI22XL U2870 ( .A0(n4137), .A1(n214), .B0(n4147), .B1(n86), .Y(n2597) );
  OAI22XL U2871 ( .A0(n4118), .A1(n470), .B0(n4127), .B1(n342), .Y(n2598) );
  OAI22XL U2872 ( .A0(n1701), .A1(n726), .B0(n1546), .B1(n598), .Y(n2595) );
  OAI22XL U2873 ( .A0(n4137), .A1(n213), .B0(n4147), .B1(n85), .Y(n2593) );
  OAI22XL U2874 ( .A0(n4118), .A1(n469), .B0(n4127), .B1(n341), .Y(n2594) );
  OAI22XL U2875 ( .A0(n1701), .A1(n725), .B0(n1546), .B1(n597), .Y(n2591) );
  OAI22XL U2876 ( .A0(n4137), .A1(n212), .B0(n4147), .B1(n84), .Y(n2589) );
  OAI22XL U2877 ( .A0(n4118), .A1(n468), .B0(n4127), .B1(n340), .Y(n2590) );
  OAI22XL U2878 ( .A0(n1701), .A1(n724), .B0(n1546), .B1(n596), .Y(n2587) );
  OAI22XL U2879 ( .A0(n4137), .A1(n211), .B0(n4147), .B1(n83), .Y(n2585) );
  OAI22XL U2880 ( .A0(n4118), .A1(n467), .B0(n4127), .B1(n339), .Y(n2586) );
  OAI22XL U2881 ( .A0(n1701), .A1(n723), .B0(n1546), .B1(n595), .Y(n2583) );
  OAI22XL U2882 ( .A0(n4137), .A1(n210), .B0(n4147), .B1(n82), .Y(n2577) );
  OAI22XL U2883 ( .A0(n4118), .A1(n466), .B0(n4127), .B1(n338), .Y(n2578) );
  OAI22XL U2884 ( .A0(n1701), .A1(n722), .B0(n1546), .B1(n594), .Y(n2575) );
  OAI22XL U2885 ( .A0(n4137), .A1(n209), .B0(n4147), .B1(n81), .Y(n2573) );
  OAI22XL U2886 ( .A0(n4118), .A1(n465), .B0(n4127), .B1(n337), .Y(n2574) );
  OAI22XL U2887 ( .A0(n1701), .A1(n721), .B0(n1546), .B1(n593), .Y(n2571) );
  OAI22XL U2888 ( .A0(n4136), .A1(n208), .B0(n4146), .B1(n80), .Y(n2569) );
  OAI22XL U2889 ( .A0(n4116), .A1(n464), .B0(n4126), .B1(n336), .Y(n2570) );
  OAI22XL U2890 ( .A0(n1558), .A1(n720), .B0(n1550), .B1(n592), .Y(n2567) );
  OAI22XL U2891 ( .A0(n4136), .A1(n207), .B0(n4146), .B1(n79), .Y(n2565) );
  OAI22XL U2892 ( .A0(n4115), .A1(n463), .B0(n4126), .B1(n335), .Y(n2566) );
  OAI22XL U2893 ( .A0(n1558), .A1(n719), .B0(n1550), .B1(n591), .Y(n2563) );
  OAI22XL U2894 ( .A0(n4136), .A1(n206), .B0(n4146), .B1(n78), .Y(n2561) );
  OAI22XL U2895 ( .A0(n4114), .A1(n462), .B0(n4126), .B1(n334), .Y(n2562) );
  OAI22XL U2896 ( .A0(n1701), .A1(n718), .B0(n1550), .B1(n590), .Y(n2559) );
  OAI22XL U2897 ( .A0(n4136), .A1(n205), .B0(n4146), .B1(n77), .Y(n2557) );
  OAI22XL U2898 ( .A0(n4112), .A1(n461), .B0(n4126), .B1(n333), .Y(n2558) );
  OAI22XL U2899 ( .A0(n1558), .A1(n717), .B0(n1546), .B1(n589), .Y(n2555) );
  OAI22XL U2900 ( .A0(n4136), .A1(n204), .B0(n4146), .B1(n76), .Y(n2553) );
  OAI22XL U2901 ( .A0(n1562), .A1(n460), .B0(n4126), .B1(n332), .Y(n2554) );
  OAI22XL U2902 ( .A0(n1696), .A1(n716), .B0(n1365), .B1(n588), .Y(n2551) );
  OAI22XL U2903 ( .A0(n4136), .A1(n203), .B0(n4146), .B1(n75), .Y(n2549) );
  OAI22XL U2904 ( .A0(n4111), .A1(n459), .B0(n4126), .B1(n331), .Y(n2550) );
  OAI22XL U2905 ( .A0(n1701), .A1(n715), .B0(n1546), .B1(n587), .Y(n2547) );
  OAI22XL U2906 ( .A0(n4136), .A1(n202), .B0(n4146), .B1(n74), .Y(n2545) );
  OAI22XL U2907 ( .A0(n1562), .A1(n458), .B0(n4126), .B1(n330), .Y(n2546) );
  OAI22XL U2908 ( .A0(n1695), .A1(n714), .B0(n1370), .B1(n586), .Y(n2543) );
  OAI22XL U2909 ( .A0(n4136), .A1(n201), .B0(n4146), .B1(n73), .Y(n2541) );
  OAI22XL U2910 ( .A0(n1562), .A1(n457), .B0(n4126), .B1(n329), .Y(n2542) );
  OAI22XL U2911 ( .A0(n1696), .A1(n713), .B0(n1358), .B1(n585), .Y(n2539) );
  OAI22XL U2912 ( .A0(n4136), .A1(n200), .B0(n4146), .B1(n72), .Y(n2533) );
  OAI22XL U2913 ( .A0(n4111), .A1(n456), .B0(n4126), .B1(n328), .Y(n2534) );
  OAI22XL U2914 ( .A0(n1701), .A1(n712), .B0(n1546), .B1(n584), .Y(n2531) );
  OAI22XL U2915 ( .A0(n4136), .A1(n199), .B0(n4146), .B1(n71), .Y(n2529) );
  OAI22XL U2916 ( .A0(n1562), .A1(n455), .B0(n4126), .B1(n327), .Y(n2530) );
  OAI22XL U2917 ( .A0(n1697), .A1(n711), .B0(n1370), .B1(n583), .Y(n2527) );
  OAI22XL U2918 ( .A0(n4136), .A1(n198), .B0(n4146), .B1(n70), .Y(n2525) );
  OAI22XL U2919 ( .A0(n4111), .A1(n454), .B0(n4126), .B1(n326), .Y(n2526) );
  OAI22XL U2920 ( .A0(n1695), .A1(n710), .B0(n1365), .B1(n582), .Y(n2523) );
  OAI22XL U2921 ( .A0(n4136), .A1(n197), .B0(n4146), .B1(n69), .Y(n2521) );
  OAI22XL U2922 ( .A0(n4111), .A1(n453), .B0(n4126), .B1(n325), .Y(n2522) );
  OAI22XL U2923 ( .A0(n1697), .A1(n709), .B0(n1528), .B1(n581), .Y(n2519) );
  OAI22XL U2924 ( .A0(n4136), .A1(n196), .B0(n4146), .B1(n68), .Y(n2517) );
  OAI22XL U2925 ( .A0(n1562), .A1(n452), .B0(n4126), .B1(n324), .Y(n2518) );
  OAI22XL U2926 ( .A0(n1701), .A1(n708), .B0(n1546), .B1(n580), .Y(n2515) );
  OAI22XL U2927 ( .A0(n4136), .A1(n195), .B0(n4146), .B1(n67), .Y(n2513) );
  OAI22XL U2928 ( .A0(n4111), .A1(n451), .B0(n4126), .B1(n323), .Y(n2514) );
  OAI22XL U2929 ( .A0(n1695), .A1(n707), .B0(n1358), .B1(n579), .Y(n2511) );
  OAI22XL U2930 ( .A0(n4136), .A1(n194), .B0(n4146), .B1(n66), .Y(n2509) );
  OAI22XL U2931 ( .A0(n1562), .A1(n450), .B0(n4126), .B1(n322), .Y(n2510) );
  OAI22XL U2932 ( .A0(n1697), .A1(n706), .B0(n1358), .B1(n578), .Y(n2507) );
  OAI22XL U2933 ( .A0(n4136), .A1(n193), .B0(n4146), .B1(n65), .Y(n2505) );
  OAI22XL U2934 ( .A0(n4111), .A1(n449), .B0(n4126), .B1(n321), .Y(n2506) );
  OAI22XL U2935 ( .A0(n1696), .A1(n705), .B0(n1370), .B1(n577), .Y(n2503) );
  OAI22XL U2936 ( .A0(n4137), .A1(n320), .B0(n4147), .B1(n192), .Y(n2625) );
  OAI22XL U2937 ( .A0(n4118), .A1(n576), .B0(n4127), .B1(n448), .Y(n2626) );
  OAI22XL U2938 ( .A0(n1701), .A1(n832), .B0(n1546), .B1(n704), .Y(n2623) );
  OAI22XL U2939 ( .A0(n4131), .A1(n319), .B0(n4145), .B1(n191), .Y(n2469) );
  OAI22XL U2940 ( .A0(n4117), .A1(n575), .B0(n1561), .B1(n447), .Y(n2470) );
  OAI22XL U2941 ( .A0(n1697), .A1(n831), .B0(n1528), .B1(n703), .Y(n2467) );
  OAI22XL U2942 ( .A0(n4134), .A1(n318), .B0(n4144), .B1(n190), .Y(n2425) );
  OAI22XL U2943 ( .A0(n4116), .A1(n574), .B0(n4124), .B1(n446), .Y(n2426) );
  OAI22XL U2944 ( .A0(n1696), .A1(n830), .B0(n1370), .B1(n702), .Y(n2423) );
  OAI22XL U2945 ( .A0(n4131), .A1(n317), .B0(n4144), .B1(n189), .Y(n2381) );
  OAI22XL U2946 ( .A0(n4116), .A1(n573), .B0(n4121), .B1(n445), .Y(n2382) );
  OAI22XL U2947 ( .A0(n1696), .A1(n829), .B0(n1370), .B1(n701), .Y(n2379) );
  OAI22XL U2948 ( .A0(n4135), .A1(n316), .B0(n4143), .B1(n188), .Y(n2337) );
  OAI22XL U2949 ( .A0(n4115), .A1(n572), .B0(n4125), .B1(n444), .Y(n2338) );
  OAI22XL U2950 ( .A0(n1695), .A1(n828), .B0(n1358), .B1(n700), .Y(n2335) );
  OAI22XL U2951 ( .A0(n4134), .A1(n315), .B0(n4142), .B1(n187), .Y(n2293) );
  OAI22XL U2952 ( .A0(n4114), .A1(n571), .B0(n4124), .B1(n443), .Y(n2294) );
  OAI22XL U2953 ( .A0(n4359), .A1(n827), .B0(n1365), .B1(n699), .Y(n2291) );
  OAI22XL U2954 ( .A0(n4136), .A1(n314), .B0(n4144), .B1(n186), .Y(n2249) );
  OAI22XL U2955 ( .A0(n4116), .A1(n570), .B0(n4126), .B1(n442), .Y(n2250) );
  OAI22XL U2956 ( .A0(n1696), .A1(n826), .B0(n1370), .B1(n698), .Y(n2247) );
  OAI22XL U2957 ( .A0(n4133), .A1(n313), .B0(n4147), .B1(n185), .Y(n2205) );
  OAI22XL U2958 ( .A0(n4113), .A1(n569), .B0(n4123), .B1(n441), .Y(n2206) );
  OAI22XL U2959 ( .A0(n1693), .A1(n825), .B0(n4357), .B1(n697), .Y(n2203) );
  OAI22XL U2960 ( .A0(n4133), .A1(n312), .B0(n4146), .B1(n184), .Y(n2161) );
  OAI22XL U2961 ( .A0(n4113), .A1(n568), .B0(n4123), .B1(n440), .Y(n2162) );
  OAI22XL U2962 ( .A0(n1693), .A1(n824), .B0(n4357), .B1(n696), .Y(n2159) );
  OAI22XL U2963 ( .A0(n4132), .A1(n311), .B0(n4141), .B1(n183), .Y(n2117) );
  OAI22XL U2964 ( .A0(n4112), .A1(n567), .B0(n4122), .B1(n439), .Y(n2118) );
  OAI22XL U2965 ( .A0(n1580), .A1(n823), .B0(n1363), .B1(n695), .Y(n2115) );
  OAI22XL U2966 ( .A0(n4137), .A1(n310), .B0(n4147), .B1(n182), .Y(n2581) );
  OAI22XL U2967 ( .A0(n4118), .A1(n566), .B0(n4127), .B1(n438), .Y(n2582) );
  OAI22XL U2968 ( .A0(n1701), .A1(n822), .B0(n1546), .B1(n694), .Y(n2579) );
  OAI22XL U2969 ( .A0(n4136), .A1(n309), .B0(n4146), .B1(n181), .Y(n2537) );
  OAI22XL U2970 ( .A0(n4116), .A1(n565), .B0(n4126), .B1(n437), .Y(n2538) );
  OAI22XL U2971 ( .A0(n4359), .A1(n821), .B0(n1550), .B1(n693), .Y(n2535) );
  OAI22XL U2972 ( .A0(n4137), .A1(n308), .B0(n4145), .B1(n180), .Y(n2501) );
  OAI22XL U2973 ( .A0(n4117), .A1(n564), .B0(n4124), .B1(n436), .Y(n2502) );
  OAI22XL U2974 ( .A0(n1697), .A1(n820), .B0(n1528), .B1(n692), .Y(n2499) );
  OAI22XL U2975 ( .A0(n4136), .A1(n307), .B0(n4145), .B1(n179), .Y(n2497) );
  OAI22XL U2976 ( .A0(n4117), .A1(n563), .B0(n4126), .B1(n435), .Y(n2498) );
  OAI22XL U2977 ( .A0(n1697), .A1(n819), .B0(n1528), .B1(n691), .Y(n2495) );
  OAI22XL U2978 ( .A0(n4134), .A1(n306), .B0(n4145), .B1(n178), .Y(n2493) );
  OAI22XL U2979 ( .A0(n4117), .A1(n562), .B0(n4122), .B1(n434), .Y(n2494) );
  OAI22XL U2980 ( .A0(n1697), .A1(n818), .B0(n1528), .B1(n690), .Y(n2491) );
  OAI22XL U2981 ( .A0(n4132), .A1(n305), .B0(n4145), .B1(n177), .Y(n2489) );
  OAI22XL U2982 ( .A0(n4117), .A1(n561), .B0(n4121), .B1(n433), .Y(n2490) );
  OAI22XL U2983 ( .A0(n1697), .A1(n817), .B0(n1528), .B1(n689), .Y(n2487) );
  OAI22XL U2984 ( .A0(n4131), .A1(n304), .B0(n4145), .B1(n176), .Y(n2485) );
  OAI22XL U2985 ( .A0(n4117), .A1(n560), .B0(n4121), .B1(n432), .Y(n2486) );
  OAI22XL U2986 ( .A0(n1697), .A1(n816), .B0(n1528), .B1(n688), .Y(n2483) );
  OAI22XL U2987 ( .A0(n4131), .A1(n303), .B0(n4145), .B1(n175), .Y(n2481) );
  OAI22XL U2988 ( .A0(n4117), .A1(n559), .B0(n4121), .B1(n431), .Y(n2482) );
  OAI22XL U2989 ( .A0(n1697), .A1(n815), .B0(n1528), .B1(n687), .Y(n2479) );
  OAI22XL U2990 ( .A0(n4135), .A1(n302), .B0(n4145), .B1(n174), .Y(n2477) );
  OAI22XL U2991 ( .A0(n4117), .A1(n558), .B0(n4127), .B1(n430), .Y(n2478) );
  OAI22XL U2992 ( .A0(n1697), .A1(n814), .B0(n1528), .B1(n686), .Y(n2475) );
  OAI22XL U2993 ( .A0(n1560), .A1(n301), .B0(n4145), .B1(n173), .Y(n2473) );
  OAI22XL U2994 ( .A0(n4117), .A1(n557), .B0(n4121), .B1(n429), .Y(n2474) );
  OAI22XL U2995 ( .A0(n1697), .A1(n813), .B0(n1528), .B1(n685), .Y(n2471) );
  OAI22XL U2996 ( .A0(n4131), .A1(n300), .B0(n4145), .B1(n172), .Y(n2465) );
  OAI22XL U2997 ( .A0(n4117), .A1(n556), .B0(n4121), .B1(n428), .Y(n2466) );
  OAI22XL U2998 ( .A0(n1697), .A1(n812), .B0(n1528), .B1(n684), .Y(n2463) );
  OAI22XL U2999 ( .A0(n4131), .A1(n299), .B0(n4145), .B1(n171), .Y(n2461) );
  OAI22XL U3000 ( .A0(n4117), .A1(n555), .B0(n4121), .B1(n427), .Y(n2462) );
  OAI22XL U3001 ( .A0(n1697), .A1(n811), .B0(n1528), .B1(n683), .Y(n2459) );
  OAI22XL U3002 ( .A0(n4131), .A1(n298), .B0(n4145), .B1(n170), .Y(n2457) );
  OAI22XL U3003 ( .A0(n4117), .A1(n554), .B0(n4121), .B1(n426), .Y(n2458) );
  OAI22XL U3004 ( .A0(n1697), .A1(n810), .B0(n1528), .B1(n682), .Y(n2455) );
  OAI22XL U3005 ( .A0(n4131), .A1(n297), .B0(n4145), .B1(n169), .Y(n2453) );
  OAI22XL U3006 ( .A0(n4117), .A1(n553), .B0(n4121), .B1(n425), .Y(n2454) );
  OAI22XL U3007 ( .A0(n1697), .A1(n809), .B0(n1528), .B1(n681), .Y(n2451) );
  OAI22XL U3008 ( .A0(n4131), .A1(n296), .B0(n4145), .B1(n168), .Y(n2449) );
  OAI22XL U3009 ( .A0(n4117), .A1(n552), .B0(n4121), .B1(n424), .Y(n2450) );
  OAI22XL U3010 ( .A0(n1697), .A1(n808), .B0(n1528), .B1(n680), .Y(n2447) );
  OAI22XL U3011 ( .A0(n4131), .A1(n295), .B0(n4145), .B1(n167), .Y(n2445) );
  OAI22XL U3012 ( .A0(n4117), .A1(n551), .B0(n4121), .B1(n423), .Y(n2446) );
  OAI22XL U3013 ( .A0(n1697), .A1(n807), .B0(n1528), .B1(n679), .Y(n2443) );
  OAI22XL U3014 ( .A0(n4131), .A1(n294), .B0(n4145), .B1(n166), .Y(n2441) );
  OAI22XL U3015 ( .A0(n4117), .A1(n550), .B0(n4121), .B1(n422), .Y(n2442) );
  OAI22XL U3016 ( .A0(n1697), .A1(n806), .B0(n1528), .B1(n678), .Y(n2439) );
  OAI22XL U3017 ( .A0(n1560), .A1(n293), .B0(n4145), .B1(n165), .Y(n2437) );
  OAI22XL U3018 ( .A0(n4117), .A1(n549), .B0(n1561), .B1(n421), .Y(n2438) );
  OAI22XL U3019 ( .A0(n1697), .A1(n805), .B0(n1528), .B1(n677), .Y(n2435) );
  OAI22XL U3020 ( .A0(n4135), .A1(n292), .B0(n4144), .B1(n164), .Y(n2433) );
  OAI22XL U3021 ( .A0(n4116), .A1(n548), .B0(n4127), .B1(n420), .Y(n2434) );
  OAI22XL U3022 ( .A0(n1696), .A1(n804), .B0(n1370), .B1(n676), .Y(n2431) );
  OAI22XL U3023 ( .A0(n4137), .A1(n291), .B0(n4144), .B1(n163), .Y(n2429) );
  OAI22XL U3024 ( .A0(n4116), .A1(n547), .B0(n4125), .B1(n419), .Y(n2430) );
  OAI22XL U3025 ( .A0(n1696), .A1(n803), .B0(n1370), .B1(n675), .Y(n2427) );
  OAI22XL U3026 ( .A0(n4136), .A1(n290), .B0(n4144), .B1(n162), .Y(n2421) );
  OAI22XL U3027 ( .A0(n4116), .A1(n546), .B0(n4126), .B1(n418), .Y(n2422) );
  OAI22XL U3028 ( .A0(n1696), .A1(n802), .B0(n1370), .B1(n674), .Y(n2419) );
  OAI22XL U3029 ( .A0(n4134), .A1(n289), .B0(n4144), .B1(n161), .Y(n2417) );
  OAI22XL U3030 ( .A0(n4116), .A1(n545), .B0(n4124), .B1(n417), .Y(n2418) );
  OAI22XL U3031 ( .A0(n1696), .A1(n801), .B0(n1370), .B1(n673), .Y(n2415) );
  OAI32X1 U3032 ( .A0(n1570), .A1(n4349), .A2(n1567), .B0(n1565), .B1(n61), 
        .Y(n3993) );
  NOR4X1 U3033 ( .A(n1571), .B(n1572), .C(n1573), .D(n1574), .Y(n1567) );
  OAI22XL U3034 ( .A0(n4132), .A1(n36), .B0(n4141), .B1(n35), .Y(n1573) );
  OAI22XL U3035 ( .A0(n1580), .A1(n40), .B0(n1363), .B1(n39), .Y(n1571) );
  OAI22XL U3036 ( .A0(n4112), .A1(n38), .B0(n4122), .B1(n37), .Y(n1574) );
  CLKBUFX3 U3037 ( .A(n4363), .Y(n1312) );
  INVXL U3038 ( .A(proc_addr[6]), .Y(n4363) );
  CLKBUFX3 U3039 ( .A(n4364), .Y(n1313) );
  INVXL U3040 ( .A(proc_addr[7]), .Y(n4364) );
  CLKBUFX3 U3041 ( .A(n4365), .Y(n1314) );
  INVXL U3042 ( .A(proc_addr[8]), .Y(n4365) );
  CLKBUFX3 U3043 ( .A(n4366), .Y(n1315) );
  INVXL U3044 ( .A(proc_addr[9]), .Y(n4366) );
  CLKBUFX3 U3045 ( .A(n4367), .Y(n1316) );
  INVXL U3046 ( .A(proc_addr[10]), .Y(n4367) );
  CLKBUFX3 U3047 ( .A(n4368), .Y(n1317) );
  INVXL U3048 ( .A(proc_addr[11]), .Y(n4368) );
  CLKBUFX3 U3049 ( .A(n4369), .Y(n1318) );
  INVXL U3050 ( .A(proc_addr[12]), .Y(n4369) );
  CLKBUFX3 U3051 ( .A(n4370), .Y(n1319) );
  INVXL U3052 ( .A(proc_addr[13]), .Y(n4370) );
  CLKBUFX3 U3053 ( .A(n4371), .Y(n1320) );
  INVXL U3054 ( .A(proc_addr[14]), .Y(n4371) );
  CLKBUFX3 U3055 ( .A(n4372), .Y(n1321) );
  INVXL U3056 ( .A(proc_addr[15]), .Y(n4372) );
  CLKBUFX3 U3057 ( .A(n4373), .Y(n1322) );
  INVXL U3058 ( .A(proc_addr[16]), .Y(n4373) );
  CLKBUFX3 U3059 ( .A(n4374), .Y(n1323) );
  INVXL U3060 ( .A(proc_addr[17]), .Y(n4374) );
  CLKBUFX3 U3061 ( .A(n4375), .Y(n1324) );
  INVXL U3062 ( .A(proc_addr[18]), .Y(n4375) );
  CLKBUFX3 U3063 ( .A(n4376), .Y(n1325) );
  INVXL U3064 ( .A(proc_addr[19]), .Y(n4376) );
  CLKBUFX3 U3065 ( .A(n4377), .Y(n1326) );
  INVXL U3066 ( .A(proc_addr[20]), .Y(n4377) );
  CLKBUFX3 U3067 ( .A(n4378), .Y(n1327) );
  INVXL U3068 ( .A(proc_addr[21]), .Y(n4378) );
  CLKBUFX3 U3069 ( .A(n4379), .Y(n1328) );
  INVXL U3070 ( .A(proc_addr[22]), .Y(n4379) );
  CLKBUFX3 U3071 ( .A(n4380), .Y(n1329) );
  INVXL U3072 ( .A(proc_addr[23]), .Y(n4380) );
  CLKBUFX3 U3073 ( .A(n4381), .Y(n1330) );
  INVXL U3074 ( .A(proc_addr[24]), .Y(n4381) );
  CLKBUFX3 U3075 ( .A(n4382), .Y(n1331) );
  INVXL U3076 ( .A(proc_addr[25]), .Y(n4382) );
  CLKBUFX3 U3077 ( .A(n4383), .Y(n1332) );
  INVXL U3078 ( .A(proc_addr[26]), .Y(n4383) );
  CLKBUFX3 U3079 ( .A(n4384), .Y(n1333) );
  INVXL U3080 ( .A(proc_addr[27]), .Y(n4384) );
  CLKBUFX3 U3081 ( .A(n4385), .Y(n1334) );
  INVXL U3082 ( .A(proc_addr[28]), .Y(n4385) );
  CLKBUFX3 U3083 ( .A(n4352), .Y(n1310) );
  INVXL U3084 ( .A(proc_addr[29]), .Y(n4352) );
  CLKBUFX3 U3085 ( .A(n4362), .Y(n1311) );
  INVXL U3086 ( .A(proc_addr[5]), .Y(n4362) );
  INVX1 U3087 ( .A(proc_wdata[18]), .Y(n4403) );
  INVX1 U3088 ( .A(proc_wdata[19]), .Y(n4404) );
  INVX1 U3089 ( .A(proc_wdata[20]), .Y(n4405) );
  INVX1 U3090 ( .A(proc_wdata[21]), .Y(n4406) );
  INVX1 U3091 ( .A(proc_wdata[22]), .Y(n4407) );
  INVX1 U3092 ( .A(proc_wdata[23]), .Y(n4408) );
  INVX1 U3093 ( .A(proc_wdata[24]), .Y(n4409) );
  INVX1 U3094 ( .A(proc_wdata[25]), .Y(n4410) );
  INVX1 U3095 ( .A(proc_wdata[26]), .Y(n4411) );
  INVX1 U3096 ( .A(proc_wdata[27]), .Y(n4412) );
  INVX1 U3097 ( .A(proc_wdata[28]), .Y(n4413) );
  INVX1 U3098 ( .A(proc_wdata[29]), .Y(n4414) );
  INVX1 U3099 ( .A(proc_wdata[30]), .Y(n4416) );
  INVX1 U3100 ( .A(proc_wdata[31]), .Y(n4415) );
  INVX1 U3101 ( .A(proc_wdata[0]), .Y(n4417) );
  INVX1 U3102 ( .A(proc_wdata[1]), .Y(n4386) );
  INVX1 U3103 ( .A(proc_wdata[2]), .Y(n4387) );
  INVX1 U3104 ( .A(proc_wdata[3]), .Y(n4388) );
  INVX1 U3105 ( .A(proc_wdata[4]), .Y(n4389) );
  INVX1 U3106 ( .A(proc_wdata[5]), .Y(n4390) );
  INVX1 U3107 ( .A(proc_wdata[6]), .Y(n4391) );
  INVX1 U3108 ( .A(proc_wdata[7]), .Y(n4392) );
  INVX1 U3109 ( .A(proc_wdata[8]), .Y(n4393) );
  INVX1 U3110 ( .A(proc_wdata[9]), .Y(n4394) );
  INVX1 U3111 ( .A(proc_wdata[10]), .Y(n4395) );
  INVX1 U3112 ( .A(proc_wdata[11]), .Y(n4396) );
  INVX1 U3113 ( .A(proc_wdata[12]), .Y(n4397) );
  INVX1 U3114 ( .A(proc_wdata[13]), .Y(n4398) );
  INVX1 U3115 ( .A(proc_wdata[14]), .Y(n4399) );
  INVX1 U3116 ( .A(proc_wdata[15]), .Y(n4400) );
  INVX1 U3117 ( .A(proc_wdata[16]), .Y(n4401) );
  INVX1 U3118 ( .A(proc_wdata[17]), .Y(n4402) );
  NOR2X1 U3119 ( .A(\state_r[0] ), .B(n4419), .Y(n1575) );
  NAND2X2 U3120 ( .A(\state_r[0] ), .B(n61), .Y(n1361) );
  NAND3X2 U3121 ( .A(n1361), .B(n61), .C(n1564), .Y(n1563) );
  NAND2X1 U3122 ( .A(n64), .B(n1576), .Y(n1564) );
  OAI22XL U3123 ( .A0(n4173), .A1(n1287), .B0(n1312), .B1(n4175), .Y(n3800) );
  OAI22XL U3124 ( .A0(n4173), .A1(n1286), .B0(n1313), .B1(n4175), .Y(n3799) );
  OAI22XL U3125 ( .A0(n4173), .A1(n1285), .B0(n1314), .B1(n4175), .Y(n3798) );
  OAI22XL U3126 ( .A0(n4173), .A1(n1284), .B0(n1315), .B1(n4176), .Y(n3797) );
  OAI22XL U3127 ( .A0(n4173), .A1(n1283), .B0(n1316), .B1(n4176), .Y(n3796) );
  OAI22XL U3128 ( .A0(n4173), .A1(n1282), .B0(n1317), .B1(n4176), .Y(n3795) );
  OAI22XL U3129 ( .A0(n4173), .A1(n1281), .B0(n1318), .B1(n4176), .Y(n3794) );
  OAI22XL U3130 ( .A0(n4173), .A1(n1280), .B0(n1319), .B1(n4175), .Y(n3793) );
  OAI22XL U3131 ( .A0(n4173), .A1(n1279), .B0(n1320), .B1(n4175), .Y(n3792) );
  OAI22XL U3132 ( .A0(n4173), .A1(n1278), .B0(n1321), .B1(n4176), .Y(n3791) );
  OAI22XL U3133 ( .A0(n4173), .A1(n1277), .B0(n1322), .B1(n4176), .Y(n3790) );
  OAI22XL U3134 ( .A0(n4174), .A1(n1276), .B0(n1323), .B1(n4176), .Y(n3789) );
  OAI22XL U3135 ( .A0(n4174), .A1(n1275), .B0(n1324), .B1(n4176), .Y(n3788) );
  OAI22XL U3136 ( .A0(n4174), .A1(n1274), .B0(n1325), .B1(n4175), .Y(n3787) );
  OAI22XL U3137 ( .A0(n4174), .A1(n1273), .B0(n1326), .B1(n4175), .Y(n3786) );
  OAI22XL U3138 ( .A0(n4174), .A1(n1272), .B0(n1327), .B1(n4175), .Y(n3785) );
  OAI22XL U3139 ( .A0(n4174), .A1(n1271), .B0(n1328), .B1(n4175), .Y(n3784) );
  OAI22XL U3140 ( .A0(n4174), .A1(n1270), .B0(n1329), .B1(n4175), .Y(n3783) );
  OAI22XL U3141 ( .A0(n4174), .A1(n1269), .B0(n1330), .B1(n4176), .Y(n3782) );
  OAI22XL U3142 ( .A0(n4174), .A1(n1268), .B0(n1331), .B1(n4175), .Y(n3781) );
  OAI22XL U3143 ( .A0(n4174), .A1(n1267), .B0(n1332), .B1(n4175), .Y(n3780) );
  OAI22XL U3144 ( .A0(n4174), .A1(n1266), .B0(n1333), .B1(n4175), .Y(n3779) );
  OAI22XL U3145 ( .A0(n4174), .A1(n1265), .B0(n1334), .B1(n4176), .Y(n3778) );
  OAI2BB2XL U3146 ( .B0(n1310), .B1(n4176), .A0N(n4176), .A1N(n1300), .Y(n3777) );
  OAI22XL U3147 ( .A0(n4149), .A1(n1113), .B0(n1311), .B1(n4152), .Y(n3975) );
  OAI22XL U3148 ( .A0(n4149), .A1(n1112), .B0(n1312), .B1(n4151), .Y(n3974) );
  OAI22XL U3149 ( .A0(n4149), .A1(n1111), .B0(n1313), .B1(n1557), .Y(n3973) );
  OAI22XL U3150 ( .A0(n4149), .A1(n1110), .B0(n1314), .B1(n4151), .Y(n3972) );
  OAI22XL U3151 ( .A0(n4149), .A1(n1109), .B0(n1315), .B1(n4152), .Y(n3971) );
  OAI22XL U3152 ( .A0(n4149), .A1(n1108), .B0(n1316), .B1(n4151), .Y(n3970) );
  OAI22XL U3153 ( .A0(n4149), .A1(n1107), .B0(n1317), .B1(n4151), .Y(n3969) );
  OAI22XL U3154 ( .A0(n4149), .A1(n1106), .B0(n1318), .B1(n4151), .Y(n3968) );
  OAI22XL U3155 ( .A0(n4149), .A1(n1105), .B0(n1319), .B1(n4151), .Y(n3967) );
  OAI22XL U3156 ( .A0(n4149), .A1(n1104), .B0(n1320), .B1(n4151), .Y(n3966) );
  OAI22XL U3157 ( .A0(n4149), .A1(n1103), .B0(n1321), .B1(n4151), .Y(n3965) );
  OAI22XL U3158 ( .A0(n4149), .A1(n1102), .B0(n1322), .B1(n4151), .Y(n3964) );
  OAI22XL U3159 ( .A0(n4150), .A1(n1101), .B0(n1323), .B1(n4152), .Y(n3963) );
  OAI22XL U3160 ( .A0(n4150), .A1(n1100), .B0(n1324), .B1(n1557), .Y(n3962) );
  OAI22XL U3161 ( .A0(n4150), .A1(n1099), .B0(n1325), .B1(n4151), .Y(n3961) );
  OAI22XL U3162 ( .A0(n4150), .A1(n1098), .B0(n1326), .B1(n4152), .Y(n3960) );
  OAI22XL U3163 ( .A0(n4150), .A1(n1097), .B0(n1327), .B1(n4152), .Y(n3959) );
  OAI22XL U3164 ( .A0(n4150), .A1(n1096), .B0(n1328), .B1(n4152), .Y(n3958) );
  OAI22XL U3165 ( .A0(n4150), .A1(n1095), .B0(n1329), .B1(n4151), .Y(n3957) );
  OAI22XL U3166 ( .A0(n4150), .A1(n1094), .B0(n1330), .B1(n4152), .Y(n3956) );
  OAI22XL U3167 ( .A0(n4150), .A1(n1093), .B0(n1331), .B1(n4152), .Y(n3955) );
  OAI22XL U3168 ( .A0(n4150), .A1(n1092), .B0(n1332), .B1(n4152), .Y(n3954) );
  OAI22XL U3169 ( .A0(n4150), .A1(n1091), .B0(n1333), .B1(n4152), .Y(n3953) );
  OAI22XL U3170 ( .A0(n4150), .A1(n1090), .B0(n1334), .B1(n4152), .Y(n3952) );
  OAI2BB2XL U3171 ( .B0(n1310), .B1(n4152), .A0N(n4151), .A1N(n1301), .Y(n3951) );
  OAI22XL U3172 ( .A0(n4153), .A1(n1138), .B0(n1311), .B1(n4155), .Y(n3950) );
  OAI22XL U3173 ( .A0(n4153), .A1(n1137), .B0(n1312), .B1(n4154), .Y(n3949) );
  OAI22XL U3174 ( .A0(n4153), .A1(n1136), .B0(n1313), .B1(n1556), .Y(n3948) );
  OAI22XL U3175 ( .A0(n4153), .A1(n1135), .B0(n1314), .B1(n4154), .Y(n3947) );
  OAI22XL U3176 ( .A0(n4153), .A1(n1134), .B0(n1315), .B1(n4155), .Y(n3946) );
  OAI22XL U3177 ( .A0(n4153), .A1(n1133), .B0(n1316), .B1(n4154), .Y(n3945) );
  OAI22XL U3178 ( .A0(n4153), .A1(n1132), .B0(n1317), .B1(n4154), .Y(n3944) );
  OAI22XL U3179 ( .A0(n4153), .A1(n1131), .B0(n1318), .B1(n4154), .Y(n3943) );
  OAI22XL U3180 ( .A0(n4153), .A1(n1130), .B0(n1319), .B1(n4154), .Y(n3942) );
  OAI22XL U3181 ( .A0(n4153), .A1(n1129), .B0(n1320), .B1(n4154), .Y(n3941) );
  OAI22XL U3182 ( .A0(n4153), .A1(n1128), .B0(n1321), .B1(n4154), .Y(n3940) );
  OAI22XL U3183 ( .A0(n4153), .A1(n1127), .B0(n1322), .B1(n4154), .Y(n3939) );
  OAI22XL U3184 ( .A0(n4153), .A1(n1126), .B0(n1323), .B1(n4155), .Y(n3938) );
  OAI22XL U3185 ( .A0(n1295), .A1(n1125), .B0(n1324), .B1(n1556), .Y(n3937) );
  OAI22XL U3186 ( .A0(n1295), .A1(n1124), .B0(n1325), .B1(n4154), .Y(n3936) );
  OAI22XL U3187 ( .A0(n4153), .A1(n1123), .B0(n1326), .B1(n4155), .Y(n3935) );
  OAI22XL U3188 ( .A0(n4153), .A1(n1122), .B0(n1327), .B1(n4155), .Y(n3934) );
  OAI22XL U3189 ( .A0(n4153), .A1(n1121), .B0(n1328), .B1(n4155), .Y(n3933) );
  OAI22XL U3190 ( .A0(n1295), .A1(n1120), .B0(n1329), .B1(n4154), .Y(n3932) );
  OAI22XL U3191 ( .A0(n4153), .A1(n1119), .B0(n1330), .B1(n4155), .Y(n3931) );
  OAI22XL U3192 ( .A0(n4153), .A1(n1118), .B0(n1331), .B1(n4155), .Y(n3930) );
  OAI22XL U3193 ( .A0(n4153), .A1(n1117), .B0(n1332), .B1(n4155), .Y(n3929) );
  OAI22XL U3194 ( .A0(n4153), .A1(n1116), .B0(n1333), .B1(n4155), .Y(n3928) );
  OAI22XL U3195 ( .A0(n4153), .A1(n1115), .B0(n1334), .B1(n4155), .Y(n3927) );
  OAI22XL U3196 ( .A0(n4156), .A1(n1163), .B0(n1311), .B1(n4158), .Y(n3925) );
  OAI22XL U3197 ( .A0(n4156), .A1(n1162), .B0(n1312), .B1(n4157), .Y(n3924) );
  OAI22XL U3198 ( .A0(n4156), .A1(n1161), .B0(n1313), .B1(n1555), .Y(n3923) );
  OAI22XL U3199 ( .A0(n4156), .A1(n1160), .B0(n1314), .B1(n4157), .Y(n3922) );
  OAI22XL U3200 ( .A0(n4156), .A1(n1159), .B0(n1315), .B1(n4158), .Y(n3921) );
  OAI22XL U3201 ( .A0(n4156), .A1(n1158), .B0(n1316), .B1(n4157), .Y(n3920) );
  OAI22XL U3202 ( .A0(n4156), .A1(n1157), .B0(n1317), .B1(n4157), .Y(n3919) );
  OAI22XL U3203 ( .A0(n4156), .A1(n1156), .B0(n1318), .B1(n4157), .Y(n3918) );
  OAI22XL U3204 ( .A0(n4156), .A1(n1155), .B0(n1319), .B1(n4157), .Y(n3917) );
  OAI22XL U3205 ( .A0(n4156), .A1(n1154), .B0(n1320), .B1(n4157), .Y(n3916) );
  OAI22XL U3206 ( .A0(n4156), .A1(n1153), .B0(n1321), .B1(n4157), .Y(n3915) );
  OAI22XL U3207 ( .A0(n4156), .A1(n1152), .B0(n1322), .B1(n4157), .Y(n3914) );
  OAI22XL U3208 ( .A0(n4156), .A1(n1151), .B0(n1323), .B1(n4158), .Y(n3913) );
  OAI22XL U3209 ( .A0(n1296), .A1(n1150), .B0(n1324), .B1(n1555), .Y(n3912) );
  OAI22XL U3210 ( .A0(n1296), .A1(n1149), .B0(n1325), .B1(n4157), .Y(n3911) );
  OAI22XL U3211 ( .A0(n4156), .A1(n1148), .B0(n1326), .B1(n4158), .Y(n3910) );
  OAI22XL U3212 ( .A0(n4156), .A1(n1147), .B0(n1327), .B1(n4158), .Y(n3909) );
  OAI22XL U3213 ( .A0(n4156), .A1(n1146), .B0(n1328), .B1(n4158), .Y(n3908) );
  OAI22XL U3214 ( .A0(n1296), .A1(n1145), .B0(n1329), .B1(n4157), .Y(n3907) );
  OAI22XL U3215 ( .A0(n4156), .A1(n1144), .B0(n1330), .B1(n4158), .Y(n3906) );
  OAI22XL U3216 ( .A0(n4156), .A1(n1143), .B0(n1331), .B1(n4158), .Y(n3905) );
  OAI22XL U3217 ( .A0(n4156), .A1(n1142), .B0(n1332), .B1(n4158), .Y(n3904) );
  OAI22XL U3218 ( .A0(n4156), .A1(n1141), .B0(n1333), .B1(n4158), .Y(n3903) );
  OAI22XL U3219 ( .A0(n4156), .A1(n1140), .B0(n1334), .B1(n4158), .Y(n3902) );
  OAI2BB2XL U3220 ( .B0(n1310), .B1(n4158), .A0N(n4157), .A1N(n1302), .Y(n3901) );
  OAI22XL U3221 ( .A0(n4159), .A1(n1188), .B0(n1311), .B1(n4160), .Y(n3900) );
  OAI22XL U3222 ( .A0(n4159), .A1(n1187), .B0(n1312), .B1(n4160), .Y(n3899) );
  OAI22XL U3223 ( .A0(n4159), .A1(n1186), .B0(n1313), .B1(n4160), .Y(n3898) );
  OAI22XL U3224 ( .A0(n4159), .A1(n1185), .B0(n1314), .B1(n4161), .Y(n3897) );
  OAI22XL U3225 ( .A0(n4159), .A1(n1184), .B0(n1315), .B1(n4161), .Y(n3896) );
  OAI22XL U3226 ( .A0(n4159), .A1(n1183), .B0(n1316), .B1(n4161), .Y(n3895) );
  OAI22XL U3227 ( .A0(n4159), .A1(n1182), .B0(n1317), .B1(n4160), .Y(n3894) );
  OAI22XL U3228 ( .A0(n4159), .A1(n1181), .B0(n1318), .B1(n1554), .Y(n3893) );
  OAI22XL U3229 ( .A0(n4159), .A1(n1180), .B0(n1319), .B1(n1554), .Y(n3892) );
  OAI22XL U3230 ( .A0(n4159), .A1(n1179), .B0(n1320), .B1(n4161), .Y(n3891) );
  OAI22XL U3231 ( .A0(n4159), .A1(n1178), .B0(n1321), .B1(n4160), .Y(n3890) );
  OAI22XL U3232 ( .A0(n4159), .A1(n1177), .B0(n1322), .B1(n4161), .Y(n3889) );
  OAI22XL U3233 ( .A0(n4159), .A1(n1176), .B0(n1323), .B1(n4161), .Y(n3888) );
  OAI22XL U3234 ( .A0(n4159), .A1(n1175), .B0(n1324), .B1(n4161), .Y(n3887) );
  OAI22XL U3235 ( .A0(n4159), .A1(n1174), .B0(n1325), .B1(n4161), .Y(n3886) );
  OAI22XL U3236 ( .A0(n4159), .A1(n1173), .B0(n1326), .B1(n4161), .Y(n3885) );
  OAI22XL U3237 ( .A0(n4159), .A1(n1172), .B0(n1327), .B1(n4161), .Y(n3884) );
  OAI22XL U3238 ( .A0(n4159), .A1(n1171), .B0(n1328), .B1(n4160), .Y(n3883) );
  OAI22XL U3239 ( .A0(n4159), .A1(n1170), .B0(n1329), .B1(n4160), .Y(n3882) );
  OAI22XL U3240 ( .A0(n4159), .A1(n1169), .B0(n1330), .B1(n4161), .Y(n3881) );
  OAI22XL U3241 ( .A0(n4159), .A1(n1168), .B0(n1331), .B1(n4160), .Y(n3880) );
  OAI22XL U3242 ( .A0(n1297), .A1(n1167), .B0(n1332), .B1(n4160), .Y(n3879) );
  OAI22XL U3243 ( .A0(n1297), .A1(n1166), .B0(n1333), .B1(n4160), .Y(n3878) );
  OAI22XL U3244 ( .A0(n1297), .A1(n1165), .B0(n1334), .B1(n4160), .Y(n3877) );
  OAI2BB2XL U3245 ( .B0(n1310), .B1(n4161), .A0N(n4160), .A1N(n1303), .Y(n3876) );
  OAI22XL U3246 ( .A0(n4162), .A1(n1213), .B0(n1311), .B1(n4164), .Y(n3875) );
  OAI22XL U3247 ( .A0(n4162), .A1(n1212), .B0(n1312), .B1(n4164), .Y(n3874) );
  OAI22XL U3248 ( .A0(n4162), .A1(n1211), .B0(n1313), .B1(n4164), .Y(n3873) );
  OAI22XL U3249 ( .A0(n4162), .A1(n1210), .B0(n1314), .B1(n4164), .Y(n3872) );
  OAI22XL U3250 ( .A0(n4162), .A1(n1209), .B0(n1315), .B1(n4165), .Y(n3871) );
  OAI22XL U3251 ( .A0(n4162), .A1(n1208), .B0(n1316), .B1(n4165), .Y(n3870) );
  OAI22XL U3252 ( .A0(n4162), .A1(n1207), .B0(n1317), .B1(n4165), .Y(n3869) );
  OAI22XL U3253 ( .A0(n4162), .A1(n1206), .B0(n1318), .B1(n4165), .Y(n3868) );
  OAI22XL U3254 ( .A0(n4162), .A1(n1205), .B0(n1319), .B1(n4164), .Y(n3867) );
  OAI22XL U3255 ( .A0(n4162), .A1(n1204), .B0(n1320), .B1(n4164), .Y(n3866) );
  OAI22XL U3256 ( .A0(n4162), .A1(n1203), .B0(n1321), .B1(n4165), .Y(n3865) );
  OAI22XL U3257 ( .A0(n4162), .A1(n1202), .B0(n1322), .B1(n4165), .Y(n3864) );
  OAI22XL U3258 ( .A0(n4163), .A1(n1201), .B0(n1323), .B1(n4165), .Y(n3863) );
  OAI22XL U3259 ( .A0(n4163), .A1(n1200), .B0(n1324), .B1(n4165), .Y(n3862) );
  OAI22XL U3260 ( .A0(n4163), .A1(n1199), .B0(n1325), .B1(n4164), .Y(n3861) );
  OAI22XL U3261 ( .A0(n4163), .A1(n1198), .B0(n1326), .B1(n4164), .Y(n3860) );
  OAI22XL U3262 ( .A0(n4163), .A1(n1197), .B0(n1327), .B1(n4164), .Y(n3859) );
  OAI22XL U3263 ( .A0(n4163), .A1(n1196), .B0(n1328), .B1(n4164), .Y(n3858) );
  OAI22XL U3264 ( .A0(n4163), .A1(n1195), .B0(n1329), .B1(n4164), .Y(n3857) );
  OAI22XL U3265 ( .A0(n4163), .A1(n1194), .B0(n1330), .B1(n4165), .Y(n3856) );
  OAI22XL U3266 ( .A0(n4163), .A1(n1193), .B0(n1331), .B1(n4164), .Y(n3855) );
  OAI22XL U3267 ( .A0(n4163), .A1(n1192), .B0(n1332), .B1(n4164), .Y(n3854) );
  OAI22XL U3268 ( .A0(n4163), .A1(n1191), .B0(n1333), .B1(n4164), .Y(n3853) );
  OAI22XL U3269 ( .A0(n4163), .A1(n1190), .B0(n1334), .B1(n4165), .Y(n3852) );
  OAI2BB2XL U3270 ( .B0(n1310), .B1(n4165), .A0N(n4165), .A1N(n1304), .Y(n3851) );
  OAI22XL U3271 ( .A0(n4166), .A1(n1238), .B0(n1311), .B1(n4168), .Y(n3850) );
  OAI22XL U3272 ( .A0(n4166), .A1(n1237), .B0(n1312), .B1(n4168), .Y(n3849) );
  OAI22XL U3273 ( .A0(n4166), .A1(n1236), .B0(n1313), .B1(n4168), .Y(n3848) );
  OAI22XL U3274 ( .A0(n4166), .A1(n1235), .B0(n1314), .B1(n4168), .Y(n3847) );
  OAI22XL U3275 ( .A0(n4166), .A1(n1234), .B0(n1315), .B1(n4169), .Y(n3846) );
  OAI22XL U3276 ( .A0(n4166), .A1(n1233), .B0(n1316), .B1(n4169), .Y(n3845) );
  OAI22XL U3277 ( .A0(n4166), .A1(n1232), .B0(n1317), .B1(n4169), .Y(n3844) );
  OAI22XL U3278 ( .A0(n4166), .A1(n1231), .B0(n1318), .B1(n4169), .Y(n3843) );
  OAI22XL U3279 ( .A0(n4166), .A1(n1230), .B0(n1319), .B1(n4168), .Y(n3842) );
  OAI22XL U3280 ( .A0(n4166), .A1(n1229), .B0(n1320), .B1(n4168), .Y(n3841) );
  OAI22XL U3281 ( .A0(n4166), .A1(n1228), .B0(n1321), .B1(n4169), .Y(n3840) );
  OAI22XL U3282 ( .A0(n4166), .A1(n1227), .B0(n1322), .B1(n4169), .Y(n3839) );
  OAI22XL U3283 ( .A0(n4167), .A1(n1226), .B0(n1323), .B1(n4169), .Y(n3838) );
  OAI22XL U3284 ( .A0(n4167), .A1(n1225), .B0(n1324), .B1(n4169), .Y(n3837) );
  OAI22XL U3285 ( .A0(n4167), .A1(n1224), .B0(n1325), .B1(n4168), .Y(n3836) );
  OAI22XL U3286 ( .A0(n4167), .A1(n1223), .B0(n1326), .B1(n4168), .Y(n3835) );
  OAI22XL U3287 ( .A0(n4167), .A1(n1222), .B0(n1327), .B1(n4168), .Y(n3834) );
  OAI22XL U3288 ( .A0(n4167), .A1(n1221), .B0(n1328), .B1(n4168), .Y(n3833) );
  OAI22XL U3289 ( .A0(n4167), .A1(n1220), .B0(n1329), .B1(n4168), .Y(n3832) );
  OAI22XL U3290 ( .A0(n4167), .A1(n1219), .B0(n1330), .B1(n4169), .Y(n3831) );
  OAI22XL U3291 ( .A0(n4167), .A1(n1218), .B0(n1331), .B1(n4168), .Y(n3830) );
  OAI22XL U3292 ( .A0(n4167), .A1(n1217), .B0(n1332), .B1(n4168), .Y(n3829) );
  OAI22XL U3293 ( .A0(n4167), .A1(n1216), .B0(n1333), .B1(n4168), .Y(n3828) );
  OAI22XL U3294 ( .A0(n4167), .A1(n1215), .B0(n1334), .B1(n4169), .Y(n3827) );
  OAI2BB2XL U3295 ( .B0(n1310), .B1(n4169), .A0N(n4169), .A1N(n1305), .Y(n3826) );
  OAI22XL U3296 ( .A0(n4170), .A1(n1263), .B0(n1311), .B1(n4172), .Y(n3825) );
  OAI22XL U3297 ( .A0(n4170), .A1(n1262), .B0(n1312), .B1(n4171), .Y(n3824) );
  OAI22XL U3298 ( .A0(n4170), .A1(n1261), .B0(n1313), .B1(n1547), .Y(n3823) );
  OAI22XL U3299 ( .A0(n4170), .A1(n1260), .B0(n1314), .B1(n4171), .Y(n3822) );
  OAI22XL U3300 ( .A0(n4170), .A1(n1259), .B0(n1315), .B1(n4172), .Y(n3821) );
  OAI22XL U3301 ( .A0(n4170), .A1(n1258), .B0(n1316), .B1(n4171), .Y(n3820) );
  OAI22XL U3302 ( .A0(n4170), .A1(n1257), .B0(n1317), .B1(n4171), .Y(n3819) );
  OAI22XL U3303 ( .A0(n4170), .A1(n1256), .B0(n1318), .B1(n4171), .Y(n3818) );
  OAI22XL U3304 ( .A0(n4170), .A1(n1255), .B0(n1319), .B1(n4171), .Y(n3817) );
  OAI22XL U3305 ( .A0(n4170), .A1(n1254), .B0(n1320), .B1(n4171), .Y(n3816) );
  OAI22XL U3306 ( .A0(n4170), .A1(n1253), .B0(n1321), .B1(n4171), .Y(n3815) );
  OAI22XL U3307 ( .A0(n4170), .A1(n1252), .B0(n1322), .B1(n4171), .Y(n3814) );
  OAI22XL U3308 ( .A0(n4170), .A1(n1251), .B0(n1323), .B1(n4172), .Y(n3813) );
  OAI22XL U3309 ( .A0(n1298), .A1(n1250), .B0(n1324), .B1(n1547), .Y(n3812) );
  OAI22XL U3310 ( .A0(n1298), .A1(n1249), .B0(n1325), .B1(n4171), .Y(n3811) );
  OAI22XL U3311 ( .A0(n4170), .A1(n1248), .B0(n1326), .B1(n4172), .Y(n3810) );
  OAI22XL U3312 ( .A0(n4170), .A1(n1247), .B0(n1327), .B1(n4172), .Y(n3809) );
  OAI22XL U3313 ( .A0(n4170), .A1(n1246), .B0(n1328), .B1(n4172), .Y(n3808) );
  OAI22XL U3314 ( .A0(n1298), .A1(n1245), .B0(n1329), .B1(n4171), .Y(n3807) );
  OAI22XL U3315 ( .A0(n4170), .A1(n1244), .B0(n1330), .B1(n4172), .Y(n3806) );
  OAI22XL U3316 ( .A0(n4170), .A1(n1243), .B0(n1331), .B1(n4172), .Y(n3805) );
  OAI22XL U3317 ( .A0(n4170), .A1(n1242), .B0(n1332), .B1(n4172), .Y(n3804) );
  OAI22XL U3318 ( .A0(n4170), .A1(n1241), .B0(n1333), .B1(n4172), .Y(n3803) );
  OAI22XL U3319 ( .A0(n4170), .A1(n1240), .B0(n1334), .B1(n4172), .Y(n3802) );
  OAI2BB2XL U3320 ( .B0(n1310), .B1(n4172), .A0N(n4171), .A1N(n1306), .Y(n3801) );
  OAI22XL U3321 ( .A0(n4173), .A1(n1288), .B0(n1311), .B1(n4175), .Y(n3994) );
  OAI21XL U3322 ( .A0(n4141), .A1(n1563), .B0(n35), .Y(n3991) );
  OAI21XL U3323 ( .A0(n4132), .A1(n1563), .B0(n36), .Y(n3990) );
  OAI21XL U3324 ( .A0(n4122), .A1(n1563), .B0(n37), .Y(n3989) );
  OAI21XL U3325 ( .A0(n4112), .A1(n1563), .B0(n38), .Y(n3988) );
  OAI21XL U3326 ( .A0(n1363), .A1(n1563), .B0(n39), .Y(n3987) );
  OAI21XL U3327 ( .A0(n1580), .A1(n1563), .B0(n40), .Y(n3986) );
  OAI21XL U3328 ( .A0(n1353), .A1(n1563), .B0(n41), .Y(n3985) );
  OAI21XL U3329 ( .A0(n2628), .A1(n1563), .B0(n42), .Y(n3984) );
  OAI21XL U3330 ( .A0(n2628), .A1(n1340), .B0(n50), .Y(n3983) );
  OAI21XL U3331 ( .A0(n1580), .A1(n1340), .B0(n48), .Y(n3981) );
  OAI21XL U3332 ( .A0(n1353), .A1(n1340), .B0(n49), .Y(n3982) );
  OAI21XL U3333 ( .A0(n1363), .A1(n1340), .B0(n47), .Y(n3980) );
  OAI21XL U3334 ( .A0(n4112), .A1(n1340), .B0(n46), .Y(n3979) );
  OAI21XL U3335 ( .A0(n4132), .A1(n1340), .B0(n44), .Y(n3977) );
  OAI21XL U3336 ( .A0(n4122), .A1(n1340), .B0(n45), .Y(n3978) );
  OAI21XL U3337 ( .A0(n4141), .A1(n1340), .B0(n43), .Y(n3976) );
  CLKINVX1 U3338 ( .A(proc_read), .Y(n4353) );
  CLKBUFX3 U3339 ( .A(n1690), .Y(n1337) );
  AOI211XL U3340 ( .A0(n4418), .A1(n1349), .B0(n4350), .C0(n4419), .Y(n1690)
         );
  CLKINVX1 U3341 ( .A(n1564), .Y(n4350) );
  CLKBUFX3 U3342 ( .A(n1559), .Y(n1340) );
  NAND3X1 U3343 ( .A(n1361), .B(n61), .C(n1568), .Y(n1559) );
  OAI2BB2XL U3344 ( .B0(n1310), .B1(n4155), .A0N(n4154), .A1N(n1307), .Y(n3926) );
  CLKINVX1 U3345 ( .A(mem_ready), .Y(n4418) );
  BUFX12 U3346 ( .A(proc_addr[3]), .Y(mem_addr[1]) );
  BUFX12 U3347 ( .A(proc_addr[2]), .Y(mem_addr[0]) );
endmodule


module cache_1 ( clk, proc_reset, proc_read, proc_write, proc_addr, proc_wdata, 
        proc_stall, proc_rdata, mem_read, mem_write, mem_addr, mem_rdata, 
        mem_wdata, mem_ready );
  input [29:0] proc_addr;
  input [31:0] proc_wdata;
  output [31:0] proc_rdata;
  output [27:0] mem_addr;
  input [127:0] mem_rdata;
  output [127:0] mem_wdata;
  input clk, proc_reset, proc_read, proc_write, mem_ready;
  output proc_stall, mem_read, mem_write;
  wire   proc_addr_1, proc_addr_0, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         \tag_r[7][18] , \tag_r[7][17] , \tag_r[7][15] , \tag_r[7][14] ,
         \tag_r[7][13] , \tag_r[7][12] , \tag_r[7][11] , \tag_r[7][6] ,
         \tag_r[7][4] , \tag_r[7][3] , \tag_r[7][2] , \tag_r[7][1] ,
         \tag_r[7][0] , \tag_r[6][18] , \tag_r[6][17] , \tag_r[6][16] ,
         \tag_r[6][15] , \tag_r[6][14] , \tag_r[6][13] , \tag_r[6][12] ,
         \tag_r[6][6] , \tag_r[6][4] , \tag_r[6][3] , \tag_r[6][2] ,
         \tag_r[6][1] , \tag_r[6][0] , \tag_r[5][18] , \tag_r[5][17] ,
         \tag_r[5][16] , \tag_r[5][15] , \tag_r[5][14] , \tag_r[5][13] ,
         \tag_r[5][12] , \tag_r[5][6] , \tag_r[5][4] , \tag_r[5][3] ,
         \tag_r[5][2] , \tag_r[5][1] , \tag_r[5][0] , \tag_r[4][18] ,
         \tag_r[4][17] , \tag_r[4][16] , \tag_r[4][15] , \tag_r[4][14] ,
         \tag_r[4][13] , \tag_r[4][12] , \tag_r[4][6] , \tag_r[4][4] ,
         \tag_r[4][3] , \tag_r[4][2] , \tag_r[4][1] , \tag_r[4][0] ,
         \tag_r[3][18] , \tag_r[3][17] , \tag_r[3][16] , \tag_r[3][15] ,
         \tag_r[3][14] , \tag_r[3][13] , \tag_r[3][12] , \tag_r[3][6] ,
         \tag_r[3][4] , \tag_r[3][3] , \tag_r[3][2] , \tag_r[3][1] ,
         \tag_r[3][0] , \tag_r[2][18] , \tag_r[2][17] , \tag_r[2][16] ,
         \tag_r[2][15] , \tag_r[2][14] , \tag_r[2][13] , \tag_r[2][12] ,
         \tag_r[2][6] , \tag_r[2][4] , \tag_r[2][3] , \tag_r[2][2] ,
         \tag_r[2][1] , \tag_r[2][0] , \tag_r[1][18] , \tag_r[1][17] ,
         \tag_r[1][16] , \tag_r[1][15] , \tag_r[1][14] , \tag_r[1][13] ,
         \tag_r[1][12] , \tag_r[1][6] , \tag_r[1][4] , \tag_r[1][3] ,
         \tag_r[1][2] , \tag_r[1][1] , \tag_r[1][0] , \tag_r[0][18] ,
         \tag_r[0][17] , \tag_r[0][15] , \tag_r[0][14] , \tag_r[0][13] ,
         \tag_r[0][12] , \tag_r[0][11] , \tag_r[0][6] , \tag_r[0][4] ,
         \tag_r[0][3] , \tag_r[0][2] , \tag_r[0][1] , \tag_r[0][0] ,
         \state_r[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n63, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1528, n1580, n1693, n1695, n1696, n1697, n1701,
         n1703, n1704, n2628, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288;
  assign proc_addr_1 = proc_addr[1];
  assign proc_addr_0 = proc_addr[0];

  DFFRX1 \dirty_r_reg[3]  ( .D(n4429), .CK(clk), .RN(n4309), .QN(n8284) );
  DFFRX1 \dirty_r_reg[2]  ( .D(n4430), .CK(clk), .RN(n4310), .QN(n8283) );
  DFFRX1 \dirty_r_reg[1]  ( .D(n4431), .CK(clk), .RN(n4310), .QN(n8282) );
  DFFRX1 \dirty_r_reg[5]  ( .D(n4427), .CK(clk), .RN(n4309), .QN(n8286) );
  DFFRX1 \dirty_r_reg[7]  ( .D(n4425), .CK(clk), .RN(n4309), .QN(n8288) );
  DFFRX1 \dirty_r_reg[0]  ( .D(n4432), .CK(clk), .RN(n4310), .QN(n8281) );
  DFFRX1 \dirty_r_reg[4]  ( .D(n4428), .CK(clk), .RN(n4309), .QN(n8285) );
  DFFRX1 \dirty_r_reg[6]  ( .D(n4426), .CK(clk), .RN(n4309), .QN(n8287) );
  DFFRX1 \block_r_reg[1][17]  ( .D(n4785), .CK(clk), .RN(n4291), .QN(n7392) );
  DFFRX1 \block_r_reg[1][16]  ( .D(n4784), .CK(clk), .RN(n4291), .QN(n7391) );
  DFFRX1 \block_r_reg[1][127]  ( .D(n4895), .CK(clk), .RN(n4279), .QN(n7502)
         );
  DFFRX1 \block_r_reg[1][126]  ( .D(n4894), .CK(clk), .RN(n4279), .QN(n7501)
         );
  DFFRX1 \block_r_reg[1][125]  ( .D(n4893), .CK(clk), .RN(n4278), .QN(n7500)
         );
  DFFRX1 \block_r_reg[1][122]  ( .D(n4890), .CK(clk), .RN(n4276), .QN(n7497)
         );
  DFFRX1 \block_r_reg[1][121]  ( .D(n4889), .CK(clk), .RN(n4275), .QN(n7496)
         );
  DFFRX1 \block_r_reg[1][120]  ( .D(n4888), .CK(clk), .RN(n4275), .QN(n7495)
         );
  DFFRX1 \block_r_reg[1][119]  ( .D(n4887), .CK(clk), .RN(n4274), .QN(n7494)
         );
  DFFRX1 \block_r_reg[1][118]  ( .D(n4886), .CK(clk), .RN(n4273), .QN(n7493)
         );
  DFFRX1 \block_r_reg[1][117]  ( .D(n4885), .CK(clk), .RN(n4273), .QN(n7492)
         );
  DFFRX1 \block_r_reg[1][116]  ( .D(n4884), .CK(clk), .RN(n4272), .QN(n7491)
         );
  DFFRX1 \block_r_reg[1][115]  ( .D(n4883), .CK(clk), .RN(n4271), .QN(n7490)
         );
  DFFRX1 \block_r_reg[1][114]  ( .D(n4882), .CK(clk), .RN(n4271), .QN(n7489)
         );
  DFFRX1 \block_r_reg[1][113]  ( .D(n4881), .CK(clk), .RN(n4270), .QN(n7488)
         );
  DFFRX1 \block_r_reg[1][112]  ( .D(n4880), .CK(clk), .RN(n4269), .QN(n7487)
         );
  DFFRX1 \block_r_reg[5][95]  ( .D(n5375), .CK(clk), .RN(n4258), .QN(n7982) );
  DFFRX1 \block_r_reg[1][95]  ( .D(n4863), .CK(clk), .RN(n4258), .QN(n7470) );
  DFFRX1 \block_r_reg[5][94]  ( .D(n5374), .CK(clk), .RN(n4258), .QN(n7981) );
  DFFRX1 \block_r_reg[1][94]  ( .D(n4862), .CK(clk), .RN(n4257), .QN(n7469) );
  DFFRX1 \block_r_reg[5][93]  ( .D(n5373), .CK(clk), .RN(n4257), .QN(n7980) );
  DFFRX1 \block_r_reg[1][93]  ( .D(n4861), .CK(clk), .RN(n4257), .QN(n7468) );
  DFFRX1 \block_r_reg[5][92]  ( .D(n5372), .CK(clk), .RN(n4256), .QN(n7979) );
  DFFRX1 \block_r_reg[1][92]  ( .D(n4860), .CK(clk), .RN(n4256), .QN(n7467) );
  DFFRX1 \block_r_reg[5][90]  ( .D(n5370), .CK(clk), .RN(n4255), .QN(n7977) );
  DFFRX1 \block_r_reg[1][90]  ( .D(n4858), .CK(clk), .RN(n4255), .QN(n7465) );
  DFFRX1 \block_r_reg[5][89]  ( .D(n5369), .CK(clk), .RN(n4254), .QN(n7976) );
  DFFRX1 \block_r_reg[1][89]  ( .D(n4857), .CK(clk), .RN(n4254), .QN(n7464) );
  DFFRX1 \block_r_reg[1][88]  ( .D(n4856), .CK(clk), .RN(n4253), .QN(n7463) );
  DFFRX1 \block_r_reg[1][87]  ( .D(n4855), .CK(clk), .RN(n4253), .QN(n7462) );
  DFFRX1 \block_r_reg[1][86]  ( .D(n4854), .CK(clk), .RN(n4252), .QN(n7461) );
  DFFRX1 \block_r_reg[1][85]  ( .D(n4853), .CK(clk), .RN(n4251), .QN(n7460) );
  DFFRX1 \block_r_reg[1][84]  ( .D(n4852), .CK(clk), .RN(n4251), .QN(n7459) );
  DFFRX1 \block_r_reg[1][83]  ( .D(n4851), .CK(clk), .RN(n4250), .QN(n7458) );
  DFFRX1 \block_r_reg[1][82]  ( .D(n4850), .CK(clk), .RN(n4249), .QN(n7457) );
  DFFRX1 \block_r_reg[1][81]  ( .D(n4849), .CK(clk), .RN(n4249), .QN(n7456) );
  DFFRX1 \block_r_reg[1][80]  ( .D(n4848), .CK(clk), .RN(n4248), .QN(n7455) );
  DFFRX1 \block_r_reg[1][63]  ( .D(n4831), .CK(clk), .RN(n4237), .QN(n7438) );
  DFFRX1 \block_r_reg[1][62]  ( .D(n4830), .CK(clk), .RN(n4236), .QN(n7437) );
  DFFRX1 \block_r_reg[1][61]  ( .D(n4829), .CK(clk), .RN(n4235), .QN(n7436) );
  DFFRX1 \block_r_reg[1][58]  ( .D(n4826), .CK(clk), .RN(n4233), .QN(n7433) );
  DFFRX1 \block_r_reg[1][57]  ( .D(n4825), .CK(clk), .RN(n4233), .QN(n7432) );
  DFFRX1 \block_r_reg[1][56]  ( .D(n4824), .CK(clk), .RN(n4232), .QN(n7431) );
  DFFRX1 \block_r_reg[1][55]  ( .D(n4823), .CK(clk), .RN(n4231), .QN(n7430) );
  DFFRX1 \block_r_reg[1][54]  ( .D(n4822), .CK(clk), .RN(n4231), .QN(n7429) );
  DFFRX1 \block_r_reg[1][53]  ( .D(n4821), .CK(clk), .RN(n4230), .QN(n7428) );
  DFFRX1 \block_r_reg[1][52]  ( .D(n4820), .CK(clk), .RN(n4229), .QN(n7427) );
  DFFRX1 \block_r_reg[1][51]  ( .D(n4819), .CK(clk), .RN(n4229), .QN(n7426) );
  DFFRX1 \block_r_reg[1][50]  ( .D(n4818), .CK(clk), .RN(n4228), .QN(n7425) );
  DFFRX1 \block_r_reg[1][49]  ( .D(n4817), .CK(clk), .RN(n4227), .QN(n7424) );
  DFFRX1 \block_r_reg[1][48]  ( .D(n4816), .CK(clk), .RN(n4227), .QN(n7423) );
  DFFRX1 \block_r_reg[1][31]  ( .D(n4799), .CK(clk), .RN(n4215), .QN(n7406) );
  DFFRX1 \block_r_reg[1][30]  ( .D(n4798), .CK(clk), .RN(n4215), .QN(n7405) );
  DFFRX1 \block_r_reg[1][29]  ( .D(n4797), .CK(clk), .RN(n4214), .QN(n7404) );
  DFFRX1 \block_r_reg[1][26]  ( .D(n4794), .CK(clk), .RN(n4212), .QN(n7401) );
  DFFRX1 \block_r_reg[1][25]  ( .D(n4793), .CK(clk), .RN(n4211), .QN(n7400) );
  DFFRX1 \block_r_reg[1][24]  ( .D(n4792), .CK(clk), .RN(n4211), .QN(n7399) );
  DFFRX1 \block_r_reg[1][23]  ( .D(n4791), .CK(clk), .RN(n4210), .QN(n7398) );
  DFFRX1 \block_r_reg[1][22]  ( .D(n4790), .CK(clk), .RN(n4209), .QN(n7397) );
  DFFRX1 \block_r_reg[1][21]  ( .D(n4789), .CK(clk), .RN(n4209), .QN(n7396) );
  DFFRX1 \block_r_reg[1][20]  ( .D(n4788), .CK(clk), .RN(n4208), .QN(n7395) );
  DFFRX1 \block_r_reg[1][19]  ( .D(n4787), .CK(clk), .RN(n4207), .QN(n7394) );
  DFFRX1 \block_r_reg[1][18]  ( .D(n4786), .CK(clk), .RN(n4207), .QN(n7393) );
  DFFRX1 \block_r_reg[7][17]  ( .D(n5553), .CK(clk), .RN(n4292), .QN(n8160) );
  DFFRX1 \block_r_reg[5][17]  ( .D(n5297), .CK(clk), .RN(n4292), .QN(n7904) );
  DFFRX1 \block_r_reg[3][17]  ( .D(n5041), .CK(clk), .RN(n4291), .QN(n7648) );
  DFFRX1 \block_r_reg[7][16]  ( .D(n5552), .CK(clk), .RN(n4291), .QN(n8159) );
  DFFRX1 \block_r_reg[5][16]  ( .D(n5296), .CK(clk), .RN(n4291), .QN(n7903) );
  DFFRX1 \block_r_reg[3][16]  ( .D(n5040), .CK(clk), .RN(n4291), .QN(n7647) );
  DFFRX1 \block_r_reg[7][127]  ( .D(n5663), .CK(clk), .RN(n4280), .QN(n8270)
         );
  DFFRX1 \block_r_reg[5][127]  ( .D(n5407), .CK(clk), .RN(n4280), .QN(n8014)
         );
  DFFRX1 \block_r_reg[4][127]  ( .D(n5279), .CK(clk), .RN(n4279), .QN(n7886)
         );
  DFFRX1 \block_r_reg[3][127]  ( .D(n5151), .CK(clk), .RN(n4279), .QN(n7758)
         );
  DFFRX1 \block_r_reg[7][126]  ( .D(n5662), .CK(clk), .RN(n4279), .QN(n8269)
         );
  DFFRX1 \block_r_reg[5][126]  ( .D(n5406), .CK(clk), .RN(n4279), .QN(n8013)
         );
  DFFRX1 \block_r_reg[4][126]  ( .D(n5278), .CK(clk), .RN(n4279), .QN(n7885)
         );
  DFFRX1 \block_r_reg[3][126]  ( .D(n5150), .CK(clk), .RN(n4279), .QN(n7757)
         );
  DFFRX1 \block_r_reg[7][125]  ( .D(n5661), .CK(clk), .RN(n4278), .QN(n8268)
         );
  DFFRX1 \block_r_reg[5][125]  ( .D(n5405), .CK(clk), .RN(n4278), .QN(n8012)
         );
  DFFRX1 \block_r_reg[4][125]  ( .D(n5277), .CK(clk), .RN(n4278), .QN(n7884)
         );
  DFFRX1 \block_r_reg[3][125]  ( .D(n5149), .CK(clk), .RN(n4278), .QN(n7756)
         );
  DFFRX1 \block_r_reg[7][122]  ( .D(n5658), .CK(clk), .RN(n4276), .QN(n8265)
         );
  DFFRX1 \block_r_reg[5][122]  ( .D(n5402), .CK(clk), .RN(n4276), .QN(n8009)
         );
  DFFRX1 \block_r_reg[4][122]  ( .D(n5274), .CK(clk), .RN(n4276), .QN(n7881)
         );
  DFFRX1 \block_r_reg[3][122]  ( .D(n5146), .CK(clk), .RN(n4276), .QN(n7753)
         );
  DFFRX1 \block_r_reg[7][121]  ( .D(n5657), .CK(clk), .RN(n4276), .QN(n8264)
         );
  DFFRX1 \block_r_reg[5][121]  ( .D(n5401), .CK(clk), .RN(n4276), .QN(n8008)
         );
  DFFRX1 \block_r_reg[4][121]  ( .D(n5273), .CK(clk), .RN(n4275), .QN(n7880)
         );
  DFFRX1 \block_r_reg[3][121]  ( .D(n5145), .CK(clk), .RN(n4275), .QN(n7752)
         );
  DFFRX1 \block_r_reg[7][120]  ( .D(n5656), .CK(clk), .RN(n4275), .QN(n8263)
         );
  DFFRX1 \block_r_reg[5][120]  ( .D(n5400), .CK(clk), .RN(n4275), .QN(n8007)
         );
  DFFRX1 \block_r_reg[4][120]  ( .D(n5272), .CK(clk), .RN(n4275), .QN(n7879)
         );
  DFFRX1 \block_r_reg[3][120]  ( .D(n5144), .CK(clk), .RN(n4275), .QN(n7751)
         );
  DFFRX1 \block_r_reg[7][119]  ( .D(n5655), .CK(clk), .RN(n4274), .QN(n8262)
         );
  DFFRX1 \block_r_reg[5][119]  ( .D(n5399), .CK(clk), .RN(n4274), .QN(n8006)
         );
  DFFRX1 \block_r_reg[4][119]  ( .D(n5271), .CK(clk), .RN(n4274), .QN(n7878)
         );
  DFFRX1 \block_r_reg[3][119]  ( .D(n5143), .CK(clk), .RN(n4274), .QN(n7750)
         );
  DFFRX1 \block_r_reg[7][118]  ( .D(n5654), .CK(clk), .RN(n4274), .QN(n8261)
         );
  DFFRX1 \block_r_reg[5][118]  ( .D(n5398), .CK(clk), .RN(n4274), .QN(n8005)
         );
  DFFRX1 \block_r_reg[4][118]  ( .D(n5270), .CK(clk), .RN(n4273), .QN(n7877)
         );
  DFFRX1 \block_r_reg[3][118]  ( .D(n5142), .CK(clk), .RN(n4273), .QN(n7749)
         );
  DFFRX1 \block_r_reg[7][117]  ( .D(n5653), .CK(clk), .RN(n4273), .QN(n8260)
         );
  DFFRX1 \block_r_reg[5][117]  ( .D(n5397), .CK(clk), .RN(n4273), .QN(n8004)
         );
  DFFRX1 \block_r_reg[3][117]  ( .D(n5141), .CK(clk), .RN(n4273), .QN(n7748)
         );
  DFFRX1 \block_r_reg[7][116]  ( .D(n5652), .CK(clk), .RN(n4272), .QN(n8259)
         );
  DFFRX1 \block_r_reg[5][116]  ( .D(n5396), .CK(clk), .RN(n4272), .QN(n8003)
         );
  DFFRX1 \block_r_reg[3][116]  ( .D(n5140), .CK(clk), .RN(n4272), .QN(n7747)
         );
  DFFRX1 \block_r_reg[7][115]  ( .D(n5651), .CK(clk), .RN(n4272), .QN(n8258)
         );
  DFFRX1 \block_r_reg[5][115]  ( .D(n5395), .CK(clk), .RN(n4272), .QN(n8002)
         );
  DFFRX1 \block_r_reg[3][115]  ( .D(n5139), .CK(clk), .RN(n4271), .QN(n7746)
         );
  DFFRX1 \block_r_reg[7][114]  ( .D(n5650), .CK(clk), .RN(n4271), .QN(n8257)
         );
  DFFRX1 \block_r_reg[5][114]  ( .D(n5394), .CK(clk), .RN(n4271), .QN(n8001)
         );
  DFFRX1 \block_r_reg[3][114]  ( .D(n5138), .CK(clk), .RN(n4271), .QN(n7745)
         );
  DFFRX1 \block_r_reg[7][113]  ( .D(n5649), .CK(clk), .RN(n4270), .QN(n8256)
         );
  DFFRX1 \block_r_reg[5][113]  ( .D(n5393), .CK(clk), .RN(n4270), .QN(n8000)
         );
  DFFRX1 \block_r_reg[3][113]  ( .D(n5137), .CK(clk), .RN(n4270), .QN(n7744)
         );
  DFFRX1 \block_r_reg[7][112]  ( .D(n5648), .CK(clk), .RN(n4270), .QN(n8255)
         );
  DFFRX1 \block_r_reg[5][112]  ( .D(n5392), .CK(clk), .RN(n4270), .QN(n7999)
         );
  DFFRX1 \block_r_reg[3][112]  ( .D(n5136), .CK(clk), .RN(n4269), .QN(n7743)
         );
  DFFRX1 \block_r_reg[7][95]  ( .D(n5631), .CK(clk), .RN(n4258), .QN(n8238) );
  DFFRX1 \block_r_reg[3][95]  ( .D(n5119), .CK(clk), .RN(n4258), .QN(n7726) );
  DFFRX1 \block_r_reg[7][94]  ( .D(n5630), .CK(clk), .RN(n4258), .QN(n8237) );
  DFFRX1 \block_r_reg[3][94]  ( .D(n5118), .CK(clk), .RN(n4257), .QN(n7725) );
  DFFRX1 \block_r_reg[7][93]  ( .D(n5629), .CK(clk), .RN(n4257), .QN(n8236) );
  DFFRX1 \block_r_reg[3][93]  ( .D(n5117), .CK(clk), .RN(n4257), .QN(n7724) );
  DFFRX1 \block_r_reg[7][92]  ( .D(n5628), .CK(clk), .RN(n4256), .QN(n8235) );
  DFFRX1 \block_r_reg[3][92]  ( .D(n5116), .CK(clk), .RN(n4256), .QN(n7723) );
  DFFRX1 \block_r_reg[7][90]  ( .D(n5626), .CK(clk), .RN(n4255), .QN(n8233) );
  DFFRX1 \block_r_reg[3][90]  ( .D(n5114), .CK(clk), .RN(n4255), .QN(n7721) );
  DFFRX1 \block_r_reg[7][89]  ( .D(n5625), .CK(clk), .RN(n4254), .QN(n8232) );
  DFFRX1 \block_r_reg[3][89]  ( .D(n5113), .CK(clk), .RN(n4254), .QN(n7720) );
  DFFRX1 \block_r_reg[7][88]  ( .D(n5624), .CK(clk), .RN(n4254), .QN(n8231) );
  DFFRX1 \block_r_reg[5][88]  ( .D(n5368), .CK(clk), .RN(n4254), .QN(n7975) );
  DFFRX1 \block_r_reg[3][88]  ( .D(n5112), .CK(clk), .RN(n4253), .QN(n7719) );
  DFFRX1 \block_r_reg[7][87]  ( .D(n5623), .CK(clk), .RN(n4253), .QN(n8230) );
  DFFRX1 \block_r_reg[5][87]  ( .D(n5367), .CK(clk), .RN(n4253), .QN(n7974) );
  DFFRX1 \block_r_reg[3][87]  ( .D(n5111), .CK(clk), .RN(n4253), .QN(n7718) );
  DFFRX1 \block_r_reg[7][86]  ( .D(n5622), .CK(clk), .RN(n4252), .QN(n8229) );
  DFFRX1 \block_r_reg[5][86]  ( .D(n5366), .CK(clk), .RN(n4252), .QN(n7973) );
  DFFRX1 \block_r_reg[3][86]  ( .D(n5110), .CK(clk), .RN(n4252), .QN(n7717) );
  DFFRX1 \block_r_reg[7][85]  ( .D(n5621), .CK(clk), .RN(n4252), .QN(n8228) );
  DFFRX1 \block_r_reg[5][85]  ( .D(n5365), .CK(clk), .RN(n4252), .QN(n7972) );
  DFFRX1 \block_r_reg[3][85]  ( .D(n5109), .CK(clk), .RN(n4251), .QN(n7716) );
  DFFRX1 \block_r_reg[7][84]  ( .D(n5620), .CK(clk), .RN(n4251), .QN(n8227) );
  DFFRX1 \block_r_reg[5][84]  ( .D(n5364), .CK(clk), .RN(n4251), .QN(n7971) );
  DFFRX1 \block_r_reg[3][84]  ( .D(n5108), .CK(clk), .RN(n4251), .QN(n7715) );
  DFFRX1 \block_r_reg[7][83]  ( .D(n5619), .CK(clk), .RN(n4250), .QN(n8226) );
  DFFRX1 \block_r_reg[5][83]  ( .D(n5363), .CK(clk), .RN(n4250), .QN(n7970) );
  DFFRX1 \block_r_reg[3][83]  ( .D(n5107), .CK(clk), .RN(n4250), .QN(n7714) );
  DFFRX1 \block_r_reg[7][82]  ( .D(n5618), .CK(clk), .RN(n4250), .QN(n8225) );
  DFFRX1 \block_r_reg[5][82]  ( .D(n5362), .CK(clk), .RN(n4250), .QN(n7969) );
  DFFRX1 \block_r_reg[3][82]  ( .D(n5106), .CK(clk), .RN(n4249), .QN(n7713) );
  DFFRX1 \block_r_reg[7][81]  ( .D(n5617), .CK(clk), .RN(n4249), .QN(n8224) );
  DFFRX1 \block_r_reg[5][81]  ( .D(n5361), .CK(clk), .RN(n4249), .QN(n7968) );
  DFFRX1 \block_r_reg[3][81]  ( .D(n5105), .CK(clk), .RN(n4249), .QN(n7712) );
  DFFRX1 \block_r_reg[7][80]  ( .D(n5616), .CK(clk), .RN(n4248), .QN(n8223) );
  DFFRX1 \block_r_reg[5][80]  ( .D(n5360), .CK(clk), .RN(n4248), .QN(n7967) );
  DFFRX1 \block_r_reg[3][80]  ( .D(n5104), .CK(clk), .RN(n4248), .QN(n7711) );
  DFFRX1 \block_r_reg[7][63]  ( .D(n5599), .CK(clk), .RN(n4237), .QN(n8206) );
  DFFRX1 \block_r_reg[5][63]  ( .D(n5343), .CK(clk), .RN(n4237), .QN(n7950) );
  DFFRX1 \block_r_reg[3][63]  ( .D(n5087), .CK(clk), .RN(n4237), .QN(n7694) );
  DFFRX1 \block_r_reg[7][62]  ( .D(n5598), .CK(clk), .RN(n4236), .QN(n8205) );
  DFFRX1 \block_r_reg[5][62]  ( .D(n5342), .CK(clk), .RN(n4236), .QN(n7949) );
  DFFRX1 \block_r_reg[3][62]  ( .D(n5086), .CK(clk), .RN(n4236), .QN(n7693) );
  DFFRX1 \block_r_reg[7][61]  ( .D(n5597), .CK(clk), .RN(n4236), .QN(n8204) );
  DFFRX1 \block_r_reg[5][61]  ( .D(n5341), .CK(clk), .RN(n4236), .QN(n7948) );
  DFFRX1 \block_r_reg[3][61]  ( .D(n5085), .CK(clk), .RN(n4235), .QN(n7692) );
  DFFRX1 \block_r_reg[7][58]  ( .D(n5594), .CK(clk), .RN(n4234), .QN(n8201) );
  DFFRX1 \block_r_reg[5][58]  ( .D(n5338), .CK(clk), .RN(n4234), .QN(n7945) );
  DFFRX1 \block_r_reg[3][58]  ( .D(n5082), .CK(clk), .RN(n4233), .QN(n7689) );
  DFFRX1 \block_r_reg[7][57]  ( .D(n5593), .CK(clk), .RN(n4233), .QN(n8200) );
  DFFRX1 \block_r_reg[5][57]  ( .D(n5337), .CK(clk), .RN(n4233), .QN(n7944) );
  DFFRX1 \block_r_reg[3][57]  ( .D(n5081), .CK(clk), .RN(n4233), .QN(n7688) );
  DFFRX1 \block_r_reg[7][56]  ( .D(n5592), .CK(clk), .RN(n4232), .QN(n8199) );
  DFFRX1 \block_r_reg[5][56]  ( .D(n5336), .CK(clk), .RN(n4232), .QN(n7943) );
  DFFRX1 \block_r_reg[3][56]  ( .D(n5080), .CK(clk), .RN(n4232), .QN(n7687) );
  DFFRX1 \block_r_reg[7][55]  ( .D(n5591), .CK(clk), .RN(n4232), .QN(n8198) );
  DFFRX1 \block_r_reg[5][55]  ( .D(n5335), .CK(clk), .RN(n4232), .QN(n7942) );
  DFFRX1 \block_r_reg[3][55]  ( .D(n5079), .CK(clk), .RN(n4231), .QN(n7686) );
  DFFRX1 \block_r_reg[7][54]  ( .D(n5590), .CK(clk), .RN(n4231), .QN(n8197) );
  DFFRX1 \block_r_reg[5][54]  ( .D(n5334), .CK(clk), .RN(n4231), .QN(n7941) );
  DFFRX1 \block_r_reg[3][54]  ( .D(n5078), .CK(clk), .RN(n4231), .QN(n7685) );
  DFFRX1 \block_r_reg[7][53]  ( .D(n5589), .CK(clk), .RN(n4230), .QN(n8196) );
  DFFRX1 \block_r_reg[5][53]  ( .D(n5333), .CK(clk), .RN(n4230), .QN(n7940) );
  DFFRX1 \block_r_reg[3][53]  ( .D(n5077), .CK(clk), .RN(n4230), .QN(n7684) );
  DFFRX1 \block_r_reg[7][52]  ( .D(n5588), .CK(clk), .RN(n4230), .QN(n8195) );
  DFFRX1 \block_r_reg[5][52]  ( .D(n5332), .CK(clk), .RN(n4230), .QN(n7939) );
  DFFRX1 \block_r_reg[3][52]  ( .D(n5076), .CK(clk), .RN(n4229), .QN(n7683) );
  DFFRX1 \block_r_reg[7][51]  ( .D(n5587), .CK(clk), .RN(n4229), .QN(n8194) );
  DFFRX1 \block_r_reg[5][51]  ( .D(n5331), .CK(clk), .RN(n4229), .QN(n7938) );
  DFFRX1 \block_r_reg[3][51]  ( .D(n5075), .CK(clk), .RN(n4229), .QN(n7682) );
  DFFRX1 \block_r_reg[7][50]  ( .D(n5586), .CK(clk), .RN(n4228), .QN(n8193) );
  DFFRX1 \block_r_reg[5][50]  ( .D(n5330), .CK(clk), .RN(n4228), .QN(n7937) );
  DFFRX1 \block_r_reg[3][50]  ( .D(n5074), .CK(clk), .RN(n4228), .QN(n7681) );
  DFFRX1 \block_r_reg[7][49]  ( .D(n5585), .CK(clk), .RN(n4228), .QN(n8192) );
  DFFRX1 \block_r_reg[5][49]  ( .D(n5329), .CK(clk), .RN(n4228), .QN(n7936) );
  DFFRX1 \block_r_reg[3][49]  ( .D(n5073), .CK(clk), .RN(n4227), .QN(n7680) );
  DFFRX1 \block_r_reg[7][48]  ( .D(n5584), .CK(clk), .RN(n4227), .QN(n8191) );
  DFFRX1 \block_r_reg[5][48]  ( .D(n5328), .CK(clk), .RN(n4227), .QN(n7935) );
  DFFRX1 \block_r_reg[3][48]  ( .D(n5072), .CK(clk), .RN(n4227), .QN(n7679) );
  DFFRX1 \block_r_reg[7][31]  ( .D(n5567), .CK(clk), .RN(n4216), .QN(n8174) );
  DFFRX1 \block_r_reg[5][31]  ( .D(n5311), .CK(clk), .RN(n4216), .QN(n7918) );
  DFFRX1 \block_r_reg[4][31]  ( .D(n5183), .CK(clk), .RN(n4215), .QN(n7790) );
  DFFRX1 \block_r_reg[3][31]  ( .D(n5055), .CK(clk), .RN(n4215), .QN(n7662) );
  DFFRX1 \block_r_reg[7][30]  ( .D(n5566), .CK(clk), .RN(n4215), .QN(n8173) );
  DFFRX1 \block_r_reg[5][30]  ( .D(n5310), .CK(clk), .RN(n4215), .QN(n7917) );
  DFFRX1 \block_r_reg[4][30]  ( .D(n5182), .CK(clk), .RN(n4215), .QN(n7789) );
  DFFRX1 \block_r_reg[3][30]  ( .D(n5054), .CK(clk), .RN(n4215), .QN(n7661) );
  DFFRX1 \block_r_reg[7][29]  ( .D(n5565), .CK(clk), .RN(n4214), .QN(n8172) );
  DFFRX1 \block_r_reg[5][29]  ( .D(n5309), .CK(clk), .RN(n4214), .QN(n7916) );
  DFFRX1 \block_r_reg[4][29]  ( .D(n5181), .CK(clk), .RN(n4214), .QN(n7788) );
  DFFRX1 \block_r_reg[3][29]  ( .D(n5053), .CK(clk), .RN(n4214), .QN(n7660) );
  DFFRX1 \block_r_reg[3][28]  ( .D(n5052), .CK(clk), .RN(n4213), .QN(n7659) );
  DFFRX1 \block_r_reg[7][26]  ( .D(n5562), .CK(clk), .RN(n4212), .QN(n8169) );
  DFFRX1 \block_r_reg[5][26]  ( .D(n5306), .CK(clk), .RN(n4212), .QN(n7913) );
  DFFRX1 \block_r_reg[4][26]  ( .D(n5178), .CK(clk), .RN(n4212), .QN(n7785) );
  DFFRX1 \block_r_reg[3][26]  ( .D(n5050), .CK(clk), .RN(n4212), .QN(n7657) );
  DFFRX1 \block_r_reg[7][25]  ( .D(n5561), .CK(clk), .RN(n4212), .QN(n8168) );
  DFFRX1 \block_r_reg[5][25]  ( .D(n5305), .CK(clk), .RN(n4212), .QN(n7912) );
  DFFRX1 \block_r_reg[4][25]  ( .D(n5177), .CK(clk), .RN(n4211), .QN(n7784) );
  DFFRX1 \block_r_reg[3][25]  ( .D(n5049), .CK(clk), .RN(n4211), .QN(n7656) );
  DFFRX1 \block_r_reg[7][24]  ( .D(n5560), .CK(clk), .RN(n4211), .QN(n8167) );
  DFFRX1 \block_r_reg[5][24]  ( .D(n5304), .CK(clk), .RN(n4211), .QN(n7911) );
  DFFRX1 \block_r_reg[4][24]  ( .D(n5176), .CK(clk), .RN(n4211), .QN(n7783) );
  DFFRX1 \block_r_reg[3][24]  ( .D(n5048), .CK(clk), .RN(n4211), .QN(n7655) );
  DFFRX1 \block_r_reg[7][23]  ( .D(n5559), .CK(clk), .RN(n4210), .QN(n8166) );
  DFFRX1 \block_r_reg[5][23]  ( .D(n5303), .CK(clk), .RN(n4210), .QN(n7910) );
  DFFRX1 \block_r_reg[4][23]  ( .D(n5175), .CK(clk), .RN(n4210), .QN(n7782) );
  DFFRX1 \block_r_reg[3][23]  ( .D(n5047), .CK(clk), .RN(n4210), .QN(n7654) );
  DFFRX1 \block_r_reg[7][22]  ( .D(n5558), .CK(clk), .RN(n4210), .QN(n8165) );
  DFFRX1 \block_r_reg[5][22]  ( .D(n5302), .CK(clk), .RN(n4210), .QN(n7909) );
  DFFRX1 \block_r_reg[4][22]  ( .D(n5174), .CK(clk), .RN(n4209), .QN(n7781) );
  DFFRX1 \block_r_reg[3][22]  ( .D(n5046), .CK(clk), .RN(n4209), .QN(n7653) );
  DFFRX1 \block_r_reg[7][21]  ( .D(n5557), .CK(clk), .RN(n4209), .QN(n8164) );
  DFFRX1 \block_r_reg[5][21]  ( .D(n5301), .CK(clk), .RN(n4209), .QN(n7908) );
  DFFRX1 \block_r_reg[4][21]  ( .D(n5173), .CK(clk), .RN(n4209), .QN(n7780) );
  DFFRX1 \block_r_reg[3][21]  ( .D(n5045), .CK(clk), .RN(n4209), .QN(n7652) );
  DFFRX1 \block_r_reg[7][20]  ( .D(n5556), .CK(clk), .RN(n4208), .QN(n8163) );
  DFFRX1 \block_r_reg[5][20]  ( .D(n5300), .CK(clk), .RN(n4208), .QN(n7907) );
  DFFRX1 \block_r_reg[4][20]  ( .D(n5172), .CK(clk), .RN(n4208), .QN(n7779) );
  DFFRX1 \block_r_reg[3][20]  ( .D(n5044), .CK(clk), .RN(n4208), .QN(n7651) );
  DFFRX1 \block_r_reg[7][19]  ( .D(n5555), .CK(clk), .RN(n4208), .QN(n8162) );
  DFFRX1 \block_r_reg[5][19]  ( .D(n5299), .CK(clk), .RN(n4208), .QN(n7906) );
  DFFRX1 \block_r_reg[4][19]  ( .D(n5171), .CK(clk), .RN(n4207), .QN(n7778) );
  DFFRX1 \block_r_reg[3][19]  ( .D(n5043), .CK(clk), .RN(n4207), .QN(n7650) );
  DFFRX1 \block_r_reg[7][18]  ( .D(n5554), .CK(clk), .RN(n4207), .QN(n8161) );
  DFFRX1 \block_r_reg[5][18]  ( .D(n5298), .CK(clk), .RN(n4207), .QN(n7905) );
  DFFRX1 \block_r_reg[3][18]  ( .D(n5042), .CK(clk), .RN(n4207), .QN(n7649) );
  DFFRX1 \block_r_reg[0][17]  ( .D(n4657), .CK(clk), .RN(n4292), .QN(n7264) );
  DFFRX1 \block_r_reg[6][17]  ( .D(n5425), .CK(clk), .RN(n4292), .QN(n8032) );
  DFFRX1 \block_r_reg[4][17]  ( .D(n5169), .CK(clk), .RN(n4291), .QN(n7776) );
  DFFRX1 \block_r_reg[2][17]  ( .D(n4913), .CK(clk), .RN(n4291), .QN(n7520) );
  DFFRX1 \block_r_reg[0][16]  ( .D(n4656), .CK(clk), .RN(n4291), .QN(n7263) );
  DFFRX1 \block_r_reg[6][16]  ( .D(n5424), .CK(clk), .RN(n4291), .QN(n8031) );
  DFFRX1 \block_r_reg[4][16]  ( .D(n5168), .CK(clk), .RN(n4291), .QN(n7775) );
  DFFRX1 \block_r_reg[2][16]  ( .D(n4912), .CK(clk), .RN(n4291), .QN(n7519) );
  DFFRX1 \block_r_reg[0][127]  ( .D(n4767), .CK(clk), .RN(n4280), .QN(n7374)
         );
  DFFRX1 \block_r_reg[6][127]  ( .D(n5535), .CK(clk), .RN(n4280), .QN(n8142)
         );
  DFFRX1 \block_r_reg[2][127]  ( .D(n5023), .CK(clk), .RN(n4279), .QN(n7630)
         );
  DFFRX1 \block_r_reg[0][126]  ( .D(n4766), .CK(clk), .RN(n4279), .QN(n7373)
         );
  DFFRX1 \block_r_reg[6][126]  ( .D(n5534), .CK(clk), .RN(n4279), .QN(n8141)
         );
  DFFRX1 \block_r_reg[2][126]  ( .D(n5022), .CK(clk), .RN(n4279), .QN(n7629)
         );
  DFFRX1 \block_r_reg[0][125]  ( .D(n4765), .CK(clk), .RN(n4278), .QN(n7372)
         );
  DFFRX1 \block_r_reg[6][125]  ( .D(n5533), .CK(clk), .RN(n4278), .QN(n8140)
         );
  DFFRX1 \block_r_reg[2][125]  ( .D(n5021), .CK(clk), .RN(n4278), .QN(n7628)
         );
  DFFRX1 \block_r_reg[2][124]  ( .D(n5020), .CK(clk), .RN(n4277), .QN(n7627)
         );
  DFFRX1 \block_r_reg[0][122]  ( .D(n4762), .CK(clk), .RN(n4276), .QN(n7369)
         );
  DFFRX1 \block_r_reg[6][122]  ( .D(n5530), .CK(clk), .RN(n4276), .QN(n8137)
         );
  DFFRX1 \block_r_reg[2][122]  ( .D(n5018), .CK(clk), .RN(n4276), .QN(n7625)
         );
  DFFRX1 \block_r_reg[0][121]  ( .D(n4761), .CK(clk), .RN(n4276), .QN(n7368)
         );
  DFFRX1 \block_r_reg[6][121]  ( .D(n5529), .CK(clk), .RN(n4276), .QN(n8136)
         );
  DFFRX1 \block_r_reg[2][121]  ( .D(n5017), .CK(clk), .RN(n4275), .QN(n7624)
         );
  DFFRX1 \block_r_reg[0][120]  ( .D(n4760), .CK(clk), .RN(n4275), .QN(n7367)
         );
  DFFRX1 \block_r_reg[6][120]  ( .D(n5528), .CK(clk), .RN(n4275), .QN(n8135)
         );
  DFFRX1 \block_r_reg[2][120]  ( .D(n5016), .CK(clk), .RN(n4275), .QN(n7623)
         );
  DFFRX1 \block_r_reg[0][119]  ( .D(n4759), .CK(clk), .RN(n4274), .QN(n7366)
         );
  DFFRX1 \block_r_reg[6][119]  ( .D(n5527), .CK(clk), .RN(n4274), .QN(n8134)
         );
  DFFRX1 \block_r_reg[2][119]  ( .D(n5015), .CK(clk), .RN(n4274), .QN(n7622)
         );
  DFFRX1 \block_r_reg[0][118]  ( .D(n4758), .CK(clk), .RN(n4274), .QN(n7365)
         );
  DFFRX1 \block_r_reg[6][118]  ( .D(n5526), .CK(clk), .RN(n4274), .QN(n8133)
         );
  DFFRX1 \block_r_reg[2][118]  ( .D(n5014), .CK(clk), .RN(n4273), .QN(n7621)
         );
  DFFRX1 \block_r_reg[0][117]  ( .D(n4757), .CK(clk), .RN(n4273), .QN(n7364)
         );
  DFFRX1 \block_r_reg[6][117]  ( .D(n5525), .CK(clk), .RN(n4273), .QN(n8132)
         );
  DFFRX1 \block_r_reg[4][117]  ( .D(n5269), .CK(clk), .RN(n4273), .QN(n7876)
         );
  DFFRX1 \block_r_reg[2][117]  ( .D(n5013), .CK(clk), .RN(n4273), .QN(n7620)
         );
  DFFRX1 \block_r_reg[0][116]  ( .D(n4756), .CK(clk), .RN(n4272), .QN(n7363)
         );
  DFFRX1 \block_r_reg[6][116]  ( .D(n5524), .CK(clk), .RN(n4272), .QN(n8131)
         );
  DFFRX1 \block_r_reg[4][116]  ( .D(n5268), .CK(clk), .RN(n4272), .QN(n7875)
         );
  DFFRX1 \block_r_reg[2][116]  ( .D(n5012), .CK(clk), .RN(n4272), .QN(n7619)
         );
  DFFRX1 \block_r_reg[0][115]  ( .D(n4755), .CK(clk), .RN(n4272), .QN(n7362)
         );
  DFFRX1 \block_r_reg[6][115]  ( .D(n5523), .CK(clk), .RN(n4272), .QN(n8130)
         );
  DFFRX1 \block_r_reg[4][115]  ( .D(n5267), .CK(clk), .RN(n4271), .QN(n7874)
         );
  DFFRX1 \block_r_reg[2][115]  ( .D(n5011), .CK(clk), .RN(n4271), .QN(n7618)
         );
  DFFRX1 \block_r_reg[0][114]  ( .D(n4754), .CK(clk), .RN(n4271), .QN(n7361)
         );
  DFFRX1 \block_r_reg[6][114]  ( .D(n5522), .CK(clk), .RN(n4271), .QN(n8129)
         );
  DFFRX1 \block_r_reg[4][114]  ( .D(n5266), .CK(clk), .RN(n4271), .QN(n7873)
         );
  DFFRX1 \block_r_reg[2][114]  ( .D(n5010), .CK(clk), .RN(n4271), .QN(n7617)
         );
  DFFRX1 \block_r_reg[0][113]  ( .D(n4753), .CK(clk), .RN(n4270), .QN(n7360)
         );
  DFFRX1 \block_r_reg[6][113]  ( .D(n5521), .CK(clk), .RN(n4270), .QN(n8128)
         );
  DFFRX1 \block_r_reg[4][113]  ( .D(n5265), .CK(clk), .RN(n4270), .QN(n7872)
         );
  DFFRX1 \block_r_reg[2][113]  ( .D(n5009), .CK(clk), .RN(n4270), .QN(n7616)
         );
  DFFRX1 \block_r_reg[0][112]  ( .D(n4752), .CK(clk), .RN(n4270), .QN(n7359)
         );
  DFFRX1 \block_r_reg[6][112]  ( .D(n5520), .CK(clk), .RN(n4270), .QN(n8127)
         );
  DFFRX1 \block_r_reg[4][112]  ( .D(n5264), .CK(clk), .RN(n4269), .QN(n7871)
         );
  DFFRX1 \block_r_reg[2][112]  ( .D(n5008), .CK(clk), .RN(n4269), .QN(n7615)
         );
  DFFRX1 \block_r_reg[0][95]  ( .D(n4735), .CK(clk), .RN(n4258), .QN(n7342) );
  DFFRX1 \block_r_reg[6][95]  ( .D(n5503), .CK(clk), .RN(n4258), .QN(n8110) );
  DFFRX1 \block_r_reg[4][95]  ( .D(n5247), .CK(clk), .RN(n4258), .QN(n7854) );
  DFFRX1 \block_r_reg[2][95]  ( .D(n4991), .CK(clk), .RN(n4258), .QN(n7598) );
  DFFRX1 \block_r_reg[0][94]  ( .D(n4734), .CK(clk), .RN(n4258), .QN(n7341) );
  DFFRX1 \block_r_reg[6][94]  ( .D(n5502), .CK(clk), .RN(n4258), .QN(n8109) );
  DFFRX1 \block_r_reg[4][94]  ( .D(n5246), .CK(clk), .RN(n4257), .QN(n7853) );
  DFFRX1 \block_r_reg[2][94]  ( .D(n4990), .CK(clk), .RN(n4257), .QN(n7597) );
  DFFRX1 \block_r_reg[0][93]  ( .D(n4733), .CK(clk), .RN(n4257), .QN(n7340) );
  DFFRX1 \block_r_reg[6][93]  ( .D(n5501), .CK(clk), .RN(n4257), .QN(n8108) );
  DFFRX1 \block_r_reg[4][93]  ( .D(n5245), .CK(clk), .RN(n4257), .QN(n7852) );
  DFFRX1 \block_r_reg[2][93]  ( .D(n4989), .CK(clk), .RN(n4257), .QN(n7596) );
  DFFRX1 \block_r_reg[0][92]  ( .D(n4732), .CK(clk), .RN(n4256), .QN(n7339) );
  DFFRX1 \block_r_reg[6][92]  ( .D(n5500), .CK(clk), .RN(n4256), .QN(n8107) );
  DFFRX1 \block_r_reg[4][92]  ( .D(n5244), .CK(clk), .RN(n4256), .QN(n7851) );
  DFFRX1 \block_r_reg[2][92]  ( .D(n4988), .CK(clk), .RN(n4256), .QN(n7595) );
  DFFRX1 \block_r_reg[0][91]  ( .D(n4731), .CK(clk), .RN(n4256), .QN(n7338) );
  DFFRX1 \block_r_reg[6][91]  ( .D(n5499), .CK(clk), .RN(n4256), .QN(n8106) );
  DFFRX1 \block_r_reg[2][91]  ( .D(n4987), .CK(clk), .RN(n4255), .QN(n7594) );
  DFFRX1 \block_r_reg[0][90]  ( .D(n4730), .CK(clk), .RN(n4255), .QN(n7337) );
  DFFRX1 \block_r_reg[6][90]  ( .D(n5498), .CK(clk), .RN(n4255), .QN(n8105) );
  DFFRX1 \block_r_reg[4][90]  ( .D(n5242), .CK(clk), .RN(n4255), .QN(n7849) );
  DFFRX1 \block_r_reg[2][90]  ( .D(n4986), .CK(clk), .RN(n4255), .QN(n7593) );
  DFFRX1 \block_r_reg[0][89]  ( .D(n4729), .CK(clk), .RN(n4254), .QN(n7336) );
  DFFRX1 \block_r_reg[6][89]  ( .D(n5497), .CK(clk), .RN(n4254), .QN(n8104) );
  DFFRX1 \block_r_reg[4][89]  ( .D(n5241), .CK(clk), .RN(n4254), .QN(n7848) );
  DFFRX1 \block_r_reg[2][89]  ( .D(n4985), .CK(clk), .RN(n4254), .QN(n7592) );
  DFFRX1 \block_r_reg[0][88]  ( .D(n4728), .CK(clk), .RN(n4254), .QN(n7335) );
  DFFRX1 \block_r_reg[6][88]  ( .D(n5496), .CK(clk), .RN(n4254), .QN(n8103) );
  DFFRX1 \block_r_reg[4][88]  ( .D(n5240), .CK(clk), .RN(n4253), .QN(n7847) );
  DFFRX1 \block_r_reg[2][88]  ( .D(n4984), .CK(clk), .RN(n4253), .QN(n7591) );
  DFFRX1 \block_r_reg[0][87]  ( .D(n4727), .CK(clk), .RN(n4253), .QN(n7334) );
  DFFRX1 \block_r_reg[6][87]  ( .D(n5495), .CK(clk), .RN(n4253), .QN(n8102) );
  DFFRX1 \block_r_reg[4][87]  ( .D(n5239), .CK(clk), .RN(n4253), .QN(n7846) );
  DFFRX1 \block_r_reg[2][87]  ( .D(n4983), .CK(clk), .RN(n4253), .QN(n7590) );
  DFFRX1 \block_r_reg[0][86]  ( .D(n4726), .CK(clk), .RN(n4252), .QN(n7333) );
  DFFRX1 \block_r_reg[6][86]  ( .D(n5494), .CK(clk), .RN(n4252), .QN(n8101) );
  DFFRX1 \block_r_reg[4][86]  ( .D(n5238), .CK(clk), .RN(n4252), .QN(n7845) );
  DFFRX1 \block_r_reg[2][86]  ( .D(n4982), .CK(clk), .RN(n4252), .QN(n7589) );
  DFFRX1 \block_r_reg[0][85]  ( .D(n4725), .CK(clk), .RN(n4252), .QN(n7332) );
  DFFRX1 \block_r_reg[6][85]  ( .D(n5493), .CK(clk), .RN(n4252), .QN(n8100) );
  DFFRX1 \block_r_reg[4][85]  ( .D(n5237), .CK(clk), .RN(n4251), .QN(n7844) );
  DFFRX1 \block_r_reg[2][85]  ( .D(n4981), .CK(clk), .RN(n4251), .QN(n7588) );
  DFFRX1 \block_r_reg[0][84]  ( .D(n4724), .CK(clk), .RN(n4251), .QN(n7331) );
  DFFRX1 \block_r_reg[6][84]  ( .D(n5492), .CK(clk), .RN(n4251), .QN(n8099) );
  DFFRX1 \block_r_reg[4][84]  ( .D(n5236), .CK(clk), .RN(n4251), .QN(n7843) );
  DFFRX1 \block_r_reg[2][84]  ( .D(n4980), .CK(clk), .RN(n4251), .QN(n7587) );
  DFFRX1 \block_r_reg[0][83]  ( .D(n4723), .CK(clk), .RN(n4250), .QN(n7330) );
  DFFRX1 \block_r_reg[6][83]  ( .D(n5491), .CK(clk), .RN(n4250), .QN(n8098) );
  DFFRX1 \block_r_reg[4][83]  ( .D(n5235), .CK(clk), .RN(n4250), .QN(n7842) );
  DFFRX1 \block_r_reg[2][83]  ( .D(n4979), .CK(clk), .RN(n4250), .QN(n7586) );
  DFFRX1 \block_r_reg[0][82]  ( .D(n4722), .CK(clk), .RN(n4250), .QN(n7329) );
  DFFRX1 \block_r_reg[6][82]  ( .D(n5490), .CK(clk), .RN(n4250), .QN(n8097) );
  DFFRX1 \block_r_reg[4][82]  ( .D(n5234), .CK(clk), .RN(n4249), .QN(n7841) );
  DFFRX1 \block_r_reg[2][82]  ( .D(n4978), .CK(clk), .RN(n4249), .QN(n7585) );
  DFFRX1 \block_r_reg[0][81]  ( .D(n4721), .CK(clk), .RN(n4249), .QN(n7328) );
  DFFRX1 \block_r_reg[6][81]  ( .D(n5489), .CK(clk), .RN(n4249), .QN(n8096) );
  DFFRX1 \block_r_reg[4][81]  ( .D(n5233), .CK(clk), .RN(n4249), .QN(n7840) );
  DFFRX1 \block_r_reg[2][81]  ( .D(n4977), .CK(clk), .RN(n4249), .QN(n7584) );
  DFFRX1 \block_r_reg[0][80]  ( .D(n4720), .CK(clk), .RN(n4248), .QN(n7327) );
  DFFRX1 \block_r_reg[6][80]  ( .D(n5488), .CK(clk), .RN(n4248), .QN(n8095) );
  DFFRX1 \block_r_reg[4][80]  ( .D(n5232), .CK(clk), .RN(n4248), .QN(n7839) );
  DFFRX1 \block_r_reg[2][80]  ( .D(n4976), .CK(clk), .RN(n4248), .QN(n7583) );
  DFFRX1 \block_r_reg[0][63]  ( .D(n4703), .CK(clk), .RN(n4237), .QN(n7310) );
  DFFRX1 \block_r_reg[6][63]  ( .D(n5471), .CK(clk), .RN(n4237), .QN(n8078) );
  DFFRX1 \block_r_reg[4][63]  ( .D(n5215), .CK(clk), .RN(n4237), .QN(n7822) );
  DFFRX1 \block_r_reg[2][63]  ( .D(n4959), .CK(clk), .RN(n4237), .QN(n7566) );
  DFFRX1 \block_r_reg[0][62]  ( .D(n4702), .CK(clk), .RN(n4236), .QN(n7309) );
  DFFRX1 \block_r_reg[6][62]  ( .D(n5470), .CK(clk), .RN(n4236), .QN(n8077) );
  DFFRX1 \block_r_reg[4][62]  ( .D(n5214), .CK(clk), .RN(n4236), .QN(n7821) );
  DFFRX1 \block_r_reg[2][62]  ( .D(n4958), .CK(clk), .RN(n4236), .QN(n7565) );
  DFFRX1 \block_r_reg[0][61]  ( .D(n4701), .CK(clk), .RN(n4236), .QN(n7308) );
  DFFRX1 \block_r_reg[6][61]  ( .D(n5469), .CK(clk), .RN(n4236), .QN(n8076) );
  DFFRX1 \block_r_reg[4][61]  ( .D(n5213), .CK(clk), .RN(n4235), .QN(n7820) );
  DFFRX1 \block_r_reg[2][61]  ( .D(n4957), .CK(clk), .RN(n4235), .QN(n7564) );
  DFFRX1 \block_r_reg[0][60]  ( .D(n4700), .CK(clk), .RN(n4235), .QN(n7307) );
  DFFRX1 \block_r_reg[6][60]  ( .D(n5468), .CK(clk), .RN(n4235), .QN(n8075) );
  DFFRX1 \block_r_reg[2][60]  ( .D(n4956), .CK(clk), .RN(n4235), .QN(n7563) );
  DFFRX1 \block_r_reg[0][58]  ( .D(n4698), .CK(clk), .RN(n4234), .QN(n7305) );
  DFFRX1 \block_r_reg[6][58]  ( .D(n5466), .CK(clk), .RN(n4234), .QN(n8073) );
  DFFRX1 \block_r_reg[4][58]  ( .D(n5210), .CK(clk), .RN(n4233), .QN(n7817) );
  DFFRX1 \block_r_reg[2][58]  ( .D(n4954), .CK(clk), .RN(n4233), .QN(n7561) );
  DFFRX1 \block_r_reg[0][57]  ( .D(n4697), .CK(clk), .RN(n4233), .QN(n7304) );
  DFFRX1 \block_r_reg[6][57]  ( .D(n5465), .CK(clk), .RN(n4233), .QN(n8072) );
  DFFRX1 \block_r_reg[4][57]  ( .D(n5209), .CK(clk), .RN(n4233), .QN(n7816) );
  DFFRX1 \block_r_reg[2][57]  ( .D(n4953), .CK(clk), .RN(n4233), .QN(n7560) );
  DFFRX1 \block_r_reg[0][56]  ( .D(n4696), .CK(clk), .RN(n4232), .QN(n7303) );
  DFFRX1 \block_r_reg[6][56]  ( .D(n5464), .CK(clk), .RN(n4232), .QN(n8071) );
  DFFRX1 \block_r_reg[4][56]  ( .D(n5208), .CK(clk), .RN(n4232), .QN(n7815) );
  DFFRX1 \block_r_reg[2][56]  ( .D(n4952), .CK(clk), .RN(n4232), .QN(n7559) );
  DFFRX1 \block_r_reg[0][55]  ( .D(n4695), .CK(clk), .RN(n4232), .QN(n7302) );
  DFFRX1 \block_r_reg[6][55]  ( .D(n5463), .CK(clk), .RN(n4232), .QN(n8070) );
  DFFRX1 \block_r_reg[4][55]  ( .D(n5207), .CK(clk), .RN(n4231), .QN(n7814) );
  DFFRX1 \block_r_reg[2][55]  ( .D(n4951), .CK(clk), .RN(n4231), .QN(n7558) );
  DFFRX1 \block_r_reg[0][54]  ( .D(n4694), .CK(clk), .RN(n4231), .QN(n7301) );
  DFFRX1 \block_r_reg[6][54]  ( .D(n5462), .CK(clk), .RN(n4231), .QN(n8069) );
  DFFRX1 \block_r_reg[4][54]  ( .D(n5206), .CK(clk), .RN(n4231), .QN(n7813) );
  DFFRX1 \block_r_reg[2][54]  ( .D(n4950), .CK(clk), .RN(n4231), .QN(n7557) );
  DFFRX1 \block_r_reg[0][53]  ( .D(n4693), .CK(clk), .RN(n4230), .QN(n7300) );
  DFFRX1 \block_r_reg[6][53]  ( .D(n5461), .CK(clk), .RN(n4230), .QN(n8068) );
  DFFRX1 \block_r_reg[4][53]  ( .D(n5205), .CK(clk), .RN(n4230), .QN(n7812) );
  DFFRX1 \block_r_reg[2][53]  ( .D(n4949), .CK(clk), .RN(n4230), .QN(n7556) );
  DFFRX1 \block_r_reg[0][52]  ( .D(n4692), .CK(clk), .RN(n4230), .QN(n7299) );
  DFFRX1 \block_r_reg[6][52]  ( .D(n5460), .CK(clk), .RN(n4230), .QN(n8067) );
  DFFRX1 \block_r_reg[4][52]  ( .D(n5204), .CK(clk), .RN(n4229), .QN(n7811) );
  DFFRX1 \block_r_reg[2][52]  ( .D(n4948), .CK(clk), .RN(n4229), .QN(n7555) );
  DFFRX1 \block_r_reg[0][51]  ( .D(n4691), .CK(clk), .RN(n4229), .QN(n7298) );
  DFFRX1 \block_r_reg[6][51]  ( .D(n5459), .CK(clk), .RN(n4229), .QN(n8066) );
  DFFRX1 \block_r_reg[4][51]  ( .D(n5203), .CK(clk), .RN(n4229), .QN(n7810) );
  DFFRX1 \block_r_reg[2][51]  ( .D(n4947), .CK(clk), .RN(n4229), .QN(n7554) );
  DFFRX1 \block_r_reg[0][50]  ( .D(n4690), .CK(clk), .RN(n4228), .QN(n7297) );
  DFFRX1 \block_r_reg[6][50]  ( .D(n5458), .CK(clk), .RN(n4228), .QN(n8065) );
  DFFRX1 \block_r_reg[4][50]  ( .D(n5202), .CK(clk), .RN(n4228), .QN(n7809) );
  DFFRX1 \block_r_reg[2][50]  ( .D(n4946), .CK(clk), .RN(n4228), .QN(n7553) );
  DFFRX1 \block_r_reg[0][49]  ( .D(n4689), .CK(clk), .RN(n4228), .QN(n7296) );
  DFFRX1 \block_r_reg[6][49]  ( .D(n5457), .CK(clk), .RN(n4228), .QN(n8064) );
  DFFRX1 \block_r_reg[4][49]  ( .D(n5201), .CK(clk), .RN(n4227), .QN(n7808) );
  DFFRX1 \block_r_reg[2][49]  ( .D(n4945), .CK(clk), .RN(n4227), .QN(n7552) );
  DFFRX1 \block_r_reg[0][48]  ( .D(n4688), .CK(clk), .RN(n4227), .QN(n7295) );
  DFFRX1 \block_r_reg[6][48]  ( .D(n5456), .CK(clk), .RN(n4227), .QN(n8063) );
  DFFRX1 \block_r_reg[4][48]  ( .D(n5200), .CK(clk), .RN(n4227), .QN(n7807) );
  DFFRX1 \block_r_reg[2][48]  ( .D(n4944), .CK(clk), .RN(n4227), .QN(n7551) );
  DFFRX1 \block_r_reg[0][31]  ( .D(n4671), .CK(clk), .RN(n4216), .QN(n7278) );
  DFFRX1 \block_r_reg[6][31]  ( .D(n5439), .CK(clk), .RN(n4216), .QN(n8046) );
  DFFRX1 \block_r_reg[2][31]  ( .D(n4927), .CK(clk), .RN(n4215), .QN(n7534) );
  DFFRX1 \block_r_reg[0][30]  ( .D(n4670), .CK(clk), .RN(n4215), .QN(n7277) );
  DFFRX1 \block_r_reg[6][30]  ( .D(n5438), .CK(clk), .RN(n4215), .QN(n8045) );
  DFFRX1 \block_r_reg[2][30]  ( .D(n4926), .CK(clk), .RN(n4215), .QN(n7533) );
  DFFRX1 \block_r_reg[0][29]  ( .D(n4669), .CK(clk), .RN(n4214), .QN(n7276) );
  DFFRX1 \block_r_reg[6][29]  ( .D(n5437), .CK(clk), .RN(n4214), .QN(n8044) );
  DFFRX1 \block_r_reg[2][29]  ( .D(n4925), .CK(clk), .RN(n4214), .QN(n7532) );
  DFFRX1 \block_r_reg[0][28]  ( .D(n4668), .CK(clk), .RN(n4214), .QN(n7275) );
  DFFRX1 \block_r_reg[2][28]  ( .D(n4924), .CK(clk), .RN(n4213), .QN(n7531) );
  DFFRX1 \block_r_reg[2][27]  ( .D(n4923), .CK(clk), .RN(n4213), .QN(n7530) );
  DFFRX1 \block_r_reg[0][26]  ( .D(n4666), .CK(clk), .RN(n4212), .QN(n7273) );
  DFFRX1 \block_r_reg[6][26]  ( .D(n5434), .CK(clk), .RN(n4212), .QN(n8041) );
  DFFRX1 \block_r_reg[2][26]  ( .D(n4922), .CK(clk), .RN(n4212), .QN(n7529) );
  DFFRX1 \block_r_reg[0][25]  ( .D(n4665), .CK(clk), .RN(n4212), .QN(n7272) );
  DFFRX1 \block_r_reg[6][25]  ( .D(n5433), .CK(clk), .RN(n4212), .QN(n8040) );
  DFFRX1 \block_r_reg[2][25]  ( .D(n4921), .CK(clk), .RN(n4211), .QN(n7528) );
  DFFRX1 \block_r_reg[0][24]  ( .D(n4664), .CK(clk), .RN(n4211), .QN(n7271) );
  DFFRX1 \block_r_reg[6][24]  ( .D(n5432), .CK(clk), .RN(n4211), .QN(n8039) );
  DFFRX1 \block_r_reg[2][24]  ( .D(n4920), .CK(clk), .RN(n4211), .QN(n7527) );
  DFFRX1 \block_r_reg[0][23]  ( .D(n4663), .CK(clk), .RN(n4210), .QN(n7270) );
  DFFRX1 \block_r_reg[6][23]  ( .D(n5431), .CK(clk), .RN(n4210), .QN(n8038) );
  DFFRX1 \block_r_reg[2][23]  ( .D(n4919), .CK(clk), .RN(n4210), .QN(n7526) );
  DFFRX1 \block_r_reg[0][22]  ( .D(n4662), .CK(clk), .RN(n4210), .QN(n7269) );
  DFFRX1 \block_r_reg[6][22]  ( .D(n5430), .CK(clk), .RN(n4210), .QN(n8037) );
  DFFRX1 \block_r_reg[2][22]  ( .D(n4918), .CK(clk), .RN(n4209), .QN(n7525) );
  DFFRX1 \block_r_reg[0][21]  ( .D(n4661), .CK(clk), .RN(n4209), .QN(n7268) );
  DFFRX1 \block_r_reg[6][21]  ( .D(n5429), .CK(clk), .RN(n4209), .QN(n8036) );
  DFFRX1 \block_r_reg[2][21]  ( .D(n4917), .CK(clk), .RN(n4209), .QN(n7524) );
  DFFRX1 \block_r_reg[0][20]  ( .D(n4660), .CK(clk), .RN(n4208), .QN(n7267) );
  DFFRX1 \block_r_reg[6][20]  ( .D(n5428), .CK(clk), .RN(n4208), .QN(n8035) );
  DFFRX1 \block_r_reg[2][20]  ( .D(n4916), .CK(clk), .RN(n4208), .QN(n7523) );
  DFFRX1 \block_r_reg[0][19]  ( .D(n4659), .CK(clk), .RN(n4208), .QN(n7266) );
  DFFRX1 \block_r_reg[6][19]  ( .D(n5427), .CK(clk), .RN(n4208), .QN(n8034) );
  DFFRX1 \block_r_reg[2][19]  ( .D(n4915), .CK(clk), .RN(n4207), .QN(n7522) );
  DFFRX1 \block_r_reg[0][18]  ( .D(n4658), .CK(clk), .RN(n4207), .QN(n7265) );
  DFFRX1 \block_r_reg[6][18]  ( .D(n5426), .CK(clk), .RN(n4207), .QN(n8033) );
  DFFRX1 \block_r_reg[4][18]  ( .D(n5170), .CK(clk), .RN(n4207), .QN(n7777) );
  DFFRX1 \block_r_reg[2][18]  ( .D(n4914), .CK(clk), .RN(n4207), .QN(n7521) );
  DFFRX1 \block_r_reg[1][124]  ( .D(n4892), .CK(clk), .RN(n4277), .QN(n7499)
         );
  DFFRX1 \block_r_reg[1][123]  ( .D(n4891), .CK(clk), .RN(n4277), .QN(n7498)
         );
  DFFRX1 \block_r_reg[5][91]  ( .D(n5371), .CK(clk), .RN(n4256), .QN(n7978) );
  DFFRX1 \block_r_reg[1][91]  ( .D(n4859), .CK(clk), .RN(n4255), .QN(n7466) );
  DFFRX1 \block_r_reg[1][60]  ( .D(n4828), .CK(clk), .RN(n4235), .QN(n7435) );
  DFFRX1 \block_r_reg[1][59]  ( .D(n4827), .CK(clk), .RN(n4234), .QN(n7434) );
  DFFRX1 \block_r_reg[1][28]  ( .D(n4796), .CK(clk), .RN(n4213), .QN(n7403) );
  DFFRX1 \block_r_reg[1][27]  ( .D(n4795), .CK(clk), .RN(n4213), .QN(n7402) );
  DFFRX1 \block_r_reg[7][124]  ( .D(n5660), .CK(clk), .RN(n4278), .QN(n8267)
         );
  DFFRX1 \block_r_reg[5][124]  ( .D(n5404), .CK(clk), .RN(n4278), .QN(n8011)
         );
  DFFRX1 \block_r_reg[4][124]  ( .D(n5276), .CK(clk), .RN(n4277), .QN(n7883)
         );
  DFFRX1 \block_r_reg[3][124]  ( .D(n5148), .CK(clk), .RN(n4277), .QN(n7755)
         );
  DFFRX1 \block_r_reg[7][123]  ( .D(n5659), .CK(clk), .RN(n4277), .QN(n8266)
         );
  DFFRX1 \block_r_reg[5][123]  ( .D(n5403), .CK(clk), .RN(n4277), .QN(n8010)
         );
  DFFRX1 \block_r_reg[4][123]  ( .D(n5275), .CK(clk), .RN(n4277), .QN(n7882)
         );
  DFFRX1 \block_r_reg[3][123]  ( .D(n5147), .CK(clk), .RN(n4277), .QN(n7754)
         );
  DFFRX1 \block_r_reg[7][91]  ( .D(n5627), .CK(clk), .RN(n4256), .QN(n8234) );
  DFFRX1 \block_r_reg[3][91]  ( .D(n5115), .CK(clk), .RN(n4255), .QN(n7722) );
  DFFRX1 \block_r_reg[7][60]  ( .D(n5596), .CK(clk), .RN(n4235), .QN(n8203) );
  DFFRX1 \block_r_reg[5][60]  ( .D(n5340), .CK(clk), .RN(n4235), .QN(n7947) );
  DFFRX1 \block_r_reg[3][60]  ( .D(n5084), .CK(clk), .RN(n4235), .QN(n7691) );
  DFFRX1 \block_r_reg[7][59]  ( .D(n5595), .CK(clk), .RN(n4234), .QN(n8202) );
  DFFRX1 \block_r_reg[5][59]  ( .D(n5339), .CK(clk), .RN(n4234), .QN(n7946) );
  DFFRX1 \block_r_reg[3][59]  ( .D(n5083), .CK(clk), .RN(n4234), .QN(n7690) );
  DFFRX1 \block_r_reg[7][28]  ( .D(n5564), .CK(clk), .RN(n4214), .QN(n8171) );
  DFFRX1 \block_r_reg[5][28]  ( .D(n5308), .CK(clk), .RN(n4214), .QN(n7915) );
  DFFRX1 \block_r_reg[4][28]  ( .D(n5180), .CK(clk), .RN(n4213), .QN(n7787) );
  DFFRX1 \block_r_reg[7][27]  ( .D(n5563), .CK(clk), .RN(n4213), .QN(n8170) );
  DFFRX1 \block_r_reg[5][27]  ( .D(n5307), .CK(clk), .RN(n4213), .QN(n7914) );
  DFFRX1 \block_r_reg[4][27]  ( .D(n5179), .CK(clk), .RN(n4213), .QN(n7786) );
  DFFRX1 \block_r_reg[3][27]  ( .D(n5051), .CK(clk), .RN(n4213), .QN(n7658) );
  DFFRX1 \block_r_reg[0][124]  ( .D(n4764), .CK(clk), .RN(n4278), .QN(n7371)
         );
  DFFRX1 \block_r_reg[6][124]  ( .D(n5532), .CK(clk), .RN(n4278), .QN(n8139)
         );
  DFFRX1 \block_r_reg[0][123]  ( .D(n4763), .CK(clk), .RN(n4277), .QN(n7370)
         );
  DFFRX1 \block_r_reg[6][123]  ( .D(n5531), .CK(clk), .RN(n4277), .QN(n8138)
         );
  DFFRX1 \block_r_reg[2][123]  ( .D(n5019), .CK(clk), .RN(n4277), .QN(n7626)
         );
  DFFRX1 \block_r_reg[4][91]  ( .D(n5243), .CK(clk), .RN(n4255), .QN(n7850) );
  DFFRX1 \block_r_reg[4][60]  ( .D(n5212), .CK(clk), .RN(n4235), .QN(n7819) );
  DFFRX1 \block_r_reg[0][59]  ( .D(n4699), .CK(clk), .RN(n4234), .QN(n7306) );
  DFFRX1 \block_r_reg[6][59]  ( .D(n5467), .CK(clk), .RN(n4234), .QN(n8074) );
  DFFRX1 \block_r_reg[4][59]  ( .D(n5211), .CK(clk), .RN(n4234), .QN(n7818) );
  DFFRX1 \block_r_reg[2][59]  ( .D(n4955), .CK(clk), .RN(n4234), .QN(n7562) );
  DFFRX1 \block_r_reg[6][28]  ( .D(n5436), .CK(clk), .RN(n4214), .QN(n8043) );
  DFFRX1 \block_r_reg[0][27]  ( .D(n4667), .CK(clk), .RN(n4213), .QN(n7274) );
  DFFRX1 \block_r_reg[6][27]  ( .D(n5435), .CK(clk), .RN(n4213), .QN(n8042) );
  DFFRX1 \valid_r_reg[7]  ( .D(n4440), .CK(clk), .RN(n4309), .QN(n8280) );
  DFFRX1 \valid_r_reg[6]  ( .D(n4439), .CK(clk), .RN(n4309), .QN(n8279) );
  DFFRX1 \valid_r_reg[5]  ( .D(n4438), .CK(clk), .RN(n4309), .QN(n8278) );
  DFFRX1 \valid_r_reg[4]  ( .D(n4437), .CK(clk), .RN(n4309), .QN(n8277) );
  DFFRX1 \valid_r_reg[3]  ( .D(n4436), .CK(clk), .RN(n4309), .QN(n8276) );
  DFFRX1 \valid_r_reg[2]  ( .D(n4435), .CK(clk), .RN(n4309), .QN(n8275) );
  DFFRX1 \valid_r_reg[1]  ( .D(n4434), .CK(clk), .RN(n4309), .QN(n8274) );
  DFFRX1 \valid_r_reg[0]  ( .D(n4433), .CK(clk), .RN(n4308), .QN(n8273) );
  DFFRX1 \tag_r_reg[3][11]  ( .D(n4552), .CK(clk), .RN(n4303), .QN(n7133) );
  DFFRX1 \tag_r_reg[3][10]  ( .D(n4551), .CK(clk), .RN(n4303), .QN(n7132) );
  DFFRX1 \tag_r_reg[3][5]  ( .D(n4546), .CK(clk), .RN(n4303), .QN(n7127) );
  DFFRX1 \tag_r_reg[7][16]  ( .D(n4457), .CK(clk), .RN(n4295), .QN(n7238) );
  DFFRX1 \tag_r_reg[7][10]  ( .D(n4451), .CK(clk), .RN(n4295), .QN(n7232) );
  DFFRX1 \tag_r_reg[7][5]  ( .D(n4446), .CK(clk), .RN(n4294), .QN(n7227) );
  DFFRX1 \tag_r_reg[2][11]  ( .D(n4577), .CK(clk), .RN(n4305), .QN(n7108) );
  DFFRX1 \tag_r_reg[2][5]  ( .D(n4571), .CK(clk), .RN(n4305), .QN(n7102) );
  DFFRX1 \tag_r_reg[0][0]  ( .D(n4422), .CK(clk), .RN(n4310), .Q(\tag_r[0][0] ), .QN(n7047) );
  DFFRX1 \tag_r_reg[1][18]  ( .D(n4609), .CK(clk), .RN(n4308), .Q(
        \tag_r[1][18] ), .QN(n7090) );
  DFFRX1 \tag_r_reg[1][17]  ( .D(n4608), .CK(clk), .RN(n4308), .Q(
        \tag_r[1][17] ), .QN(n7089) );
  DFFRX1 \tag_r_reg[1][16]  ( .D(n4607), .CK(clk), .RN(n4308), .Q(
        \tag_r[1][16] ), .QN(n7088) );
  DFFRX1 \tag_r_reg[1][15]  ( .D(n4606), .CK(clk), .RN(n4308), .Q(
        \tag_r[1][15] ), .QN(n7087) );
  DFFRX1 \tag_r_reg[1][14]  ( .D(n4605), .CK(clk), .RN(n4308), .Q(
        \tag_r[1][14] ), .QN(n7086) );
  DFFRX1 \tag_r_reg[1][13]  ( .D(n4604), .CK(clk), .RN(n4307), .Q(
        \tag_r[1][13] ), .QN(n7085) );
  DFFRX1 \tag_r_reg[1][12]  ( .D(n4603), .CK(clk), .RN(n4307), .Q(
        \tag_r[1][12] ), .QN(n7084) );
  DFFRX1 \tag_r_reg[1][6]  ( .D(n4597), .CK(clk), .RN(n4307), .Q(\tag_r[1][6] ), .QN(n7078) );
  DFFRX1 \tag_r_reg[1][4]  ( .D(n4595), .CK(clk), .RN(n4307), .Q(\tag_r[1][4] ), .QN(n7076) );
  DFFRX1 \tag_r_reg[1][3]  ( .D(n4594), .CK(clk), .RN(n4307), .Q(\tag_r[1][3] ), .QN(n7075) );
  DFFRX1 \tag_r_reg[1][2]  ( .D(n4593), .CK(clk), .RN(n4307), .Q(\tag_r[1][2] ), .QN(n7074) );
  DFFRX1 \tag_r_reg[1][1]  ( .D(n4592), .CK(clk), .RN(n4306), .Q(\tag_r[1][1] ), .QN(n7073) );
  DFFRX1 \tag_r_reg[1][0]  ( .D(n4591), .CK(clk), .RN(n4306), .Q(\tag_r[1][0] ), .QN(n7072) );
  DFFRX1 \tag_r_reg[2][18]  ( .D(n4584), .CK(clk), .RN(n4306), .Q(
        \tag_r[2][18] ), .QN(n7115) );
  DFFRX1 \tag_r_reg[2][17]  ( .D(n4583), .CK(clk), .RN(n4306), .Q(
        \tag_r[2][17] ), .QN(n7114) );
  DFFRX1 \tag_r_reg[2][16]  ( .D(n4582), .CK(clk), .RN(n4306), .Q(
        \tag_r[2][16] ), .QN(n7113) );
  DFFRX1 \tag_r_reg[2][15]  ( .D(n4581), .CK(clk), .RN(n4306), .Q(
        \tag_r[2][15] ), .QN(n7112) );
  DFFRX1 \tag_r_reg[2][14]  ( .D(n4580), .CK(clk), .RN(n4305), .Q(
        \tag_r[2][14] ), .QN(n7111) );
  DFFRX1 \tag_r_reg[2][13]  ( .D(n4579), .CK(clk), .RN(n4305), .Q(
        \tag_r[2][13] ), .QN(n7110) );
  DFFRX1 \tag_r_reg[2][12]  ( .D(n4578), .CK(clk), .RN(n4305), .Q(
        \tag_r[2][12] ), .QN(n7109) );
  DFFRX1 \tag_r_reg[2][6]  ( .D(n4572), .CK(clk), .RN(n4305), .Q(\tag_r[2][6] ), .QN(n7103) );
  DFFRX1 \tag_r_reg[2][4]  ( .D(n4570), .CK(clk), .RN(n4305), .Q(\tag_r[2][4] ), .QN(n7101) );
  DFFRX1 \tag_r_reg[2][3]  ( .D(n4569), .CK(clk), .RN(n4305), .Q(\tag_r[2][3] ), .QN(n7100) );
  DFFRX1 \tag_r_reg[2][2]  ( .D(n4568), .CK(clk), .RN(n4304), .Q(\tag_r[2][2] ), .QN(n7099) );
  DFFRX1 \tag_r_reg[2][1]  ( .D(n4567), .CK(clk), .RN(n4304), .Q(\tag_r[2][1] ), .QN(n7098) );
  DFFRX1 \tag_r_reg[2][0]  ( .D(n4566), .CK(clk), .RN(n4304), .Q(\tag_r[2][0] ), .QN(n7097) );
  DFFRX1 \tag_r_reg[3][18]  ( .D(n4559), .CK(clk), .RN(n4304), .Q(
        \tag_r[3][18] ), .QN(n7140) );
  DFFRX1 \tag_r_reg[3][17]  ( .D(n4558), .CK(clk), .RN(n4304), .Q(
        \tag_r[3][17] ), .QN(n7139) );
  DFFRX1 \tag_r_reg[3][16]  ( .D(n4557), .CK(clk), .RN(n4304), .Q(
        \tag_r[3][16] ), .QN(n7138) );
  DFFRX1 \tag_r_reg[3][15]  ( .D(n4556), .CK(clk), .RN(n4303), .Q(
        \tag_r[3][15] ), .QN(n7137) );
  DFFRX1 \tag_r_reg[3][14]  ( .D(n4555), .CK(clk), .RN(n4303), .Q(
        \tag_r[3][14] ), .QN(n7136) );
  DFFRX1 \tag_r_reg[3][13]  ( .D(n4554), .CK(clk), .RN(n4303), .Q(
        \tag_r[3][13] ), .QN(n7135) );
  DFFRX1 \tag_r_reg[3][12]  ( .D(n4553), .CK(clk), .RN(n4303), .Q(
        \tag_r[3][12] ), .QN(n7134) );
  DFFRX1 \tag_r_reg[3][6]  ( .D(n4547), .CK(clk), .RN(n4303), .Q(\tag_r[3][6] ), .QN(n7128) );
  DFFRX1 \tag_r_reg[3][4]  ( .D(n4545), .CK(clk), .RN(n4303), .Q(\tag_r[3][4] ), .QN(n7126) );
  DFFRX1 \tag_r_reg[3][3]  ( .D(n4544), .CK(clk), .RN(n4302), .Q(\tag_r[3][3] ), .QN(n7125) );
  DFFRX1 \tag_r_reg[3][2]  ( .D(n4543), .CK(clk), .RN(n4302), .Q(\tag_r[3][2] ), .QN(n7124) );
  DFFRX1 \tag_r_reg[3][1]  ( .D(n4542), .CK(clk), .RN(n4302), .Q(\tag_r[3][1] ), .QN(n7123) );
  DFFRX1 \tag_r_reg[3][0]  ( .D(n4541), .CK(clk), .RN(n4302), .Q(\tag_r[3][0] ), .QN(n7122) );
  DFFRX1 \tag_r_reg[4][18]  ( .D(n4534), .CK(clk), .RN(n4302), .Q(
        \tag_r[4][18] ), .QN(n7165) );
  DFFRX1 \tag_r_reg[4][17]  ( .D(n4533), .CK(clk), .RN(n4302), .Q(
        \tag_r[4][17] ), .QN(n7164) );
  DFFRX1 \tag_r_reg[4][16]  ( .D(n4532), .CK(clk), .RN(n4301), .Q(
        \tag_r[4][16] ), .QN(n7163) );
  DFFRX1 \tag_r_reg[4][15]  ( .D(n4531), .CK(clk), .RN(n4301), .Q(
        \tag_r[4][15] ), .QN(n7162) );
  DFFRX1 \tag_r_reg[4][14]  ( .D(n4530), .CK(clk), .RN(n4301), .Q(
        \tag_r[4][14] ), .QN(n7161) );
  DFFRX1 \tag_r_reg[4][13]  ( .D(n4529), .CK(clk), .RN(n4301), .Q(
        \tag_r[4][13] ), .QN(n7160) );
  DFFRX1 \tag_r_reg[4][12]  ( .D(n4528), .CK(clk), .RN(n4301), .Q(
        \tag_r[4][12] ), .QN(n7159) );
  DFFRX1 \tag_r_reg[4][6]  ( .D(n4522), .CK(clk), .RN(n4301), .Q(\tag_r[4][6] ), .QN(n7153) );
  DFFRX1 \tag_r_reg[4][4]  ( .D(n4520), .CK(clk), .RN(n4300), .Q(\tag_r[4][4] ), .QN(n7151) );
  DFFRX1 \tag_r_reg[4][3]  ( .D(n4519), .CK(clk), .RN(n4300), .Q(\tag_r[4][3] ), .QN(n7150) );
  DFFRX1 \tag_r_reg[4][2]  ( .D(n4518), .CK(clk), .RN(n4300), .Q(\tag_r[4][2] ), .QN(n7149) );
  DFFRX1 \tag_r_reg[4][1]  ( .D(n4517), .CK(clk), .RN(n4300), .Q(\tag_r[4][1] ), .QN(n7148) );
  DFFRX1 \tag_r_reg[4][0]  ( .D(n4516), .CK(clk), .RN(n4300), .Q(\tag_r[4][0] ), .QN(n7147) );
  DFFRX1 \tag_r_reg[5][18]  ( .D(n4509), .CK(clk), .RN(n4300), .Q(
        \tag_r[5][18] ), .QN(n7190) );
  DFFRX1 \tag_r_reg[5][17]  ( .D(n4508), .CK(clk), .RN(n4299), .Q(
        \tag_r[5][17] ), .QN(n7189) );
  DFFRX1 \tag_r_reg[5][16]  ( .D(n4507), .CK(clk), .RN(n4299), .Q(
        \tag_r[5][16] ), .QN(n7188) );
  DFFRX1 \tag_r_reg[5][15]  ( .D(n4506), .CK(clk), .RN(n4299), .Q(
        \tag_r[5][15] ), .QN(n7187) );
  DFFRX1 \tag_r_reg[5][14]  ( .D(n4505), .CK(clk), .RN(n4299), .Q(
        \tag_r[5][14] ), .QN(n7186) );
  DFFRX1 \tag_r_reg[5][13]  ( .D(n4504), .CK(clk), .RN(n4299), .Q(
        \tag_r[5][13] ), .QN(n7185) );
  DFFRX1 \tag_r_reg[5][12]  ( .D(n4503), .CK(clk), .RN(n4299), .Q(
        \tag_r[5][12] ), .QN(n7184) );
  DFFRX1 \tag_r_reg[5][6]  ( .D(n4497), .CK(clk), .RN(n4299), .Q(\tag_r[5][6] ), .QN(n7178) );
  DFFRX1 \tag_r_reg[5][4]  ( .D(n4495), .CK(clk), .RN(n4298), .Q(\tag_r[5][4] ), .QN(n7176) );
  DFFRX1 \tag_r_reg[5][3]  ( .D(n4494), .CK(clk), .RN(n4298), .Q(\tag_r[5][3] ), .QN(n7175) );
  DFFRX1 \tag_r_reg[5][2]  ( .D(n4493), .CK(clk), .RN(n4298), .Q(\tag_r[5][2] ), .QN(n7174) );
  DFFRX1 \tag_r_reg[5][1]  ( .D(n4492), .CK(clk), .RN(n4298), .Q(\tag_r[5][1] ), .QN(n7173) );
  DFFRX1 \tag_r_reg[5][0]  ( .D(n4491), .CK(clk), .RN(n4298), .Q(\tag_r[5][0] ), .QN(n7172) );
  DFFRX1 \tag_r_reg[6][18]  ( .D(n4484), .CK(clk), .RN(n4297), .Q(
        \tag_r[6][18] ), .QN(n7215) );
  DFFRX1 \tag_r_reg[6][17]  ( .D(n4483), .CK(clk), .RN(n4297), .Q(
        \tag_r[6][17] ), .QN(n7214) );
  DFFRX1 \tag_r_reg[6][16]  ( .D(n4482), .CK(clk), .RN(n4297), .Q(
        \tag_r[6][16] ), .QN(n7213) );
  DFFRX1 \tag_r_reg[6][15]  ( .D(n4481), .CK(clk), .RN(n4297), .Q(
        \tag_r[6][15] ), .QN(n7212) );
  DFFRX1 \tag_r_reg[6][14]  ( .D(n4480), .CK(clk), .RN(n4297), .Q(
        \tag_r[6][14] ), .QN(n7211) );
  DFFRX1 \tag_r_reg[6][13]  ( .D(n4479), .CK(clk), .RN(n4297), .Q(
        \tag_r[6][13] ), .QN(n7210) );
  DFFRX1 \tag_r_reg[6][12]  ( .D(n4478), .CK(clk), .RN(n4297), .Q(
        \tag_r[6][12] ), .QN(n7209) );
  DFFRX1 \tag_r_reg[6][6]  ( .D(n4472), .CK(clk), .RN(n4296), .Q(\tag_r[6][6] ), .QN(n7203) );
  DFFRX1 \tag_r_reg[6][4]  ( .D(n4470), .CK(clk), .RN(n4296), .Q(\tag_r[6][4] ), .QN(n7201) );
  DFFRX1 \tag_r_reg[6][3]  ( .D(n4469), .CK(clk), .RN(n4296), .Q(\tag_r[6][3] ), .QN(n7200) );
  DFFRX1 \tag_r_reg[6][2]  ( .D(n4468), .CK(clk), .RN(n4296), .Q(\tag_r[6][2] ), .QN(n7199) );
  DFFRX1 \tag_r_reg[6][1]  ( .D(n4467), .CK(clk), .RN(n4296), .Q(\tag_r[6][1] ), .QN(n7198) );
  DFFRX1 \tag_r_reg[6][0]  ( .D(n4466), .CK(clk), .RN(n4296), .Q(\tag_r[6][0] ), .QN(n7197) );
  DFFRX1 \tag_r_reg[7][18]  ( .D(n4459), .CK(clk), .RN(n4295), .Q(
        \tag_r[7][18] ), .QN(n7240) );
  DFFRX1 \tag_r_reg[7][17]  ( .D(n4458), .CK(clk), .RN(n4295), .Q(
        \tag_r[7][17] ), .QN(n7239) );
  DFFRX1 \tag_r_reg[7][15]  ( .D(n4456), .CK(clk), .RN(n4295), .Q(
        \tag_r[7][15] ), .QN(n7237) );
  DFFRX1 \tag_r_reg[7][14]  ( .D(n4455), .CK(clk), .RN(n4295), .Q(
        \tag_r[7][14] ), .QN(n7236) );
  DFFRX1 \tag_r_reg[7][13]  ( .D(n4454), .CK(clk), .RN(n4295), .Q(
        \tag_r[7][13] ), .QN(n7235) );
  DFFRX1 \tag_r_reg[7][12]  ( .D(n4453), .CK(clk), .RN(n4295), .Q(
        \tag_r[7][12] ), .QN(n7234) );
  DFFRX1 \tag_r_reg[7][11]  ( .D(n4452), .CK(clk), .RN(n4295), .Q(
        \tag_r[7][11] ), .QN(n7233) );
  DFFRX1 \tag_r_reg[7][6]  ( .D(n4447), .CK(clk), .RN(n4294), .Q(\tag_r[7][6] ), .QN(n7228) );
  DFFRX1 \tag_r_reg[7][4]  ( .D(n4445), .CK(clk), .RN(n4294), .Q(\tag_r[7][4] ), .QN(n7226) );
  DFFRX1 \tag_r_reg[7][3]  ( .D(n4444), .CK(clk), .RN(n4294), .Q(\tag_r[7][3] ), .QN(n7225) );
  DFFRX1 \tag_r_reg[7][2]  ( .D(n4443), .CK(clk), .RN(n4294), .Q(\tag_r[7][2] ), .QN(n7224) );
  DFFRX1 \tag_r_reg[7][1]  ( .D(n4442), .CK(clk), .RN(n4294), .Q(\tag_r[7][1] ), .QN(n7223) );
  DFFRX1 \tag_r_reg[7][0]  ( .D(n4441), .CK(clk), .RN(n4294), .Q(\tag_r[7][0] ), .QN(n7222) );
  DFFRX1 \tag_r_reg[0][18]  ( .D(n4633), .CK(clk), .RN(n4293), .Q(
        \tag_r[0][18] ), .QN(n7065) );
  DFFRX1 \tag_r_reg[0][17]  ( .D(n4632), .CK(clk), .RN(n4293), .Q(
        \tag_r[0][17] ), .QN(n7064) );
  DFFRX1 \tag_r_reg[0][15]  ( .D(n4630), .CK(clk), .RN(n4293), .Q(
        \tag_r[0][15] ), .QN(n7062) );
  DFFRX1 \tag_r_reg[0][14]  ( .D(n4629), .CK(clk), .RN(n4293), .Q(
        \tag_r[0][14] ), .QN(n7061) );
  DFFRX1 \tag_r_reg[0][13]  ( .D(n4628), .CK(clk), .RN(n4293), .Q(
        \tag_r[0][13] ), .QN(n7060) );
  DFFRX1 \tag_r_reg[0][12]  ( .D(n4627), .CK(clk), .RN(n4293), .Q(
        \tag_r[0][12] ), .QN(n7059) );
  DFFRX1 \tag_r_reg[0][11]  ( .D(n4626), .CK(clk), .RN(n4293), .Q(
        \tag_r[0][11] ), .QN(n7058) );
  DFFRX1 \tag_r_reg[0][6]  ( .D(n4621), .CK(clk), .RN(n4292), .Q(\tag_r[0][6] ), .QN(n7053) );
  DFFRX1 \tag_r_reg[0][4]  ( .D(n4619), .CK(clk), .RN(n4292), .Q(\tag_r[0][4] ), .QN(n7051) );
  DFFRX1 \tag_r_reg[0][3]  ( .D(n4618), .CK(clk), .RN(n4292), .Q(\tag_r[0][3] ), .QN(n7050) );
  DFFRX1 \tag_r_reg[0][2]  ( .D(n4617), .CK(clk), .RN(n4292), .Q(\tag_r[0][2] ), .QN(n7049) );
  DFFRX1 \tag_r_reg[0][1]  ( .D(n4616), .CK(clk), .RN(n4292), .Q(\tag_r[0][1] ), .QN(n7048) );
  DFFRX1 \block_r_reg[1][15]  ( .D(n4783), .CK(clk), .RN(n4290), .QN(n7390) );
  DFFRX1 \block_r_reg[1][14]  ( .D(n4782), .CK(clk), .RN(n4289), .QN(n7389) );
  DFFRX1 \block_r_reg[1][13]  ( .D(n4781), .CK(clk), .RN(n4289), .QN(n7388) );
  DFFRX1 \block_r_reg[1][12]  ( .D(n4780), .CK(clk), .RN(n4288), .QN(n7387) );
  DFFRX1 \block_r_reg[1][11]  ( .D(n4779), .CK(clk), .RN(n4287), .QN(n7386) );
  DFFRX1 \block_r_reg[1][10]  ( .D(n4778), .CK(clk), .RN(n4287), .QN(n7385) );
  DFFRX1 \block_r_reg[1][9]  ( .D(n4777), .CK(clk), .RN(n4286), .QN(n7384) );
  DFFRX1 \block_r_reg[1][111]  ( .D(n4879), .CK(clk), .RN(n4269), .QN(n7486)
         );
  DFFRX1 \block_r_reg[1][110]  ( .D(n4878), .CK(clk), .RN(n4268), .QN(n7485)
         );
  DFFRX1 \block_r_reg[1][109]  ( .D(n4877), .CK(clk), .RN(n4267), .QN(n7484)
         );
  DFFRX1 \block_r_reg[1][108]  ( .D(n4876), .CK(clk), .RN(n4267), .QN(n7483)
         );
  DFFRX1 \block_r_reg[1][107]  ( .D(n4875), .CK(clk), .RN(n4266), .QN(n7482)
         );
  DFFRX1 \block_r_reg[1][106]  ( .D(n4874), .CK(clk), .RN(n4265), .QN(n7481)
         );
  DFFRX1 \block_r_reg[1][105]  ( .D(n4873), .CK(clk), .RN(n4265), .QN(n7480)
         );
  DFFRX1 \block_r_reg[1][79]  ( .D(n4847), .CK(clk), .RN(n4247), .QN(n7454) );
  DFFRX1 \block_r_reg[1][78]  ( .D(n4846), .CK(clk), .RN(n4247), .QN(n7453) );
  DFFRX1 \block_r_reg[1][77]  ( .D(n4845), .CK(clk), .RN(n4246), .QN(n7452) );
  DFFRX1 \block_r_reg[1][76]  ( .D(n4844), .CK(clk), .RN(n4245), .QN(n7451) );
  DFFRX1 \block_r_reg[1][75]  ( .D(n4843), .CK(clk), .RN(n4245), .QN(n7450) );
  DFFRX1 \block_r_reg[1][74]  ( .D(n4842), .CK(clk), .RN(n4244), .QN(n7449) );
  DFFRX1 \block_r_reg[1][73]  ( .D(n4841), .CK(clk), .RN(n4243), .QN(n7448) );
  DFFRX1 \block_r_reg[1][72]  ( .D(n4840), .CK(clk), .RN(n4243), .QN(n7447) );
  DFFRX1 \block_r_reg[1][47]  ( .D(n4815), .CK(clk), .RN(n4226), .QN(n7422) );
  DFFRX1 \block_r_reg[1][46]  ( .D(n4814), .CK(clk), .RN(n4225), .QN(n7421) );
  DFFRX1 \block_r_reg[1][45]  ( .D(n4813), .CK(clk), .RN(n4225), .QN(n7420) );
  DFFRX1 \block_r_reg[1][44]  ( .D(n4812), .CK(clk), .RN(n4224), .QN(n7419) );
  DFFRX1 \block_r_reg[1][43]  ( .D(n4811), .CK(clk), .RN(n4223), .QN(n7418) );
  DFFRX1 \block_r_reg[1][42]  ( .D(n4810), .CK(clk), .RN(n4223), .QN(n7417) );
  DFFRX1 \block_r_reg[1][41]  ( .D(n4809), .CK(clk), .RN(n4222), .QN(n7416) );
  DFFRX1 \block_r_reg[1][40]  ( .D(n4808), .CK(clk), .RN(n4221), .QN(n7415) );
  DFFRX1 \block_r_reg[7][15]  ( .D(n5551), .CK(clk), .RN(n4290), .QN(n8158) );
  DFFRX1 \block_r_reg[5][15]  ( .D(n5295), .CK(clk), .RN(n4290), .QN(n7902) );
  DFFRX1 \block_r_reg[3][15]  ( .D(n5039), .CK(clk), .RN(n4290), .QN(n7646) );
  DFFRX1 \block_r_reg[7][14]  ( .D(n5550), .CK(clk), .RN(n4290), .QN(n8157) );
  DFFRX1 \block_r_reg[5][14]  ( .D(n5294), .CK(clk), .RN(n4290), .QN(n7901) );
  DFFRX1 \block_r_reg[3][14]  ( .D(n5038), .CK(clk), .RN(n4289), .QN(n7645) );
  DFFRX1 \block_r_reg[7][13]  ( .D(n5549), .CK(clk), .RN(n4289), .QN(n8156) );
  DFFRX1 \block_r_reg[5][13]  ( .D(n5293), .CK(clk), .RN(n4289), .QN(n7900) );
  DFFRX1 \block_r_reg[3][13]  ( .D(n5037), .CK(clk), .RN(n4289), .QN(n7644) );
  DFFRX1 \block_r_reg[7][12]  ( .D(n5548), .CK(clk), .RN(n4288), .QN(n8155) );
  DFFRX1 \block_r_reg[5][12]  ( .D(n5292), .CK(clk), .RN(n4288), .QN(n7899) );
  DFFRX1 \block_r_reg[3][12]  ( .D(n5036), .CK(clk), .RN(n4288), .QN(n7643) );
  DFFRX1 \block_r_reg[7][11]  ( .D(n5547), .CK(clk), .RN(n4288), .QN(n8154) );
  DFFRX1 \block_r_reg[5][11]  ( .D(n5291), .CK(clk), .RN(n4288), .QN(n7898) );
  DFFRX1 \block_r_reg[3][11]  ( .D(n5035), .CK(clk), .RN(n4287), .QN(n7642) );
  DFFRX1 \block_r_reg[7][10]  ( .D(n5546), .CK(clk), .RN(n4287), .QN(n8153) );
  DFFRX1 \block_r_reg[5][10]  ( .D(n5290), .CK(clk), .RN(n4287), .QN(n7897) );
  DFFRX1 \block_r_reg[3][10]  ( .D(n5034), .CK(clk), .RN(n4287), .QN(n7641) );
  DFFRX1 \block_r_reg[7][9]  ( .D(n5545), .CK(clk), .RN(n4286), .QN(n8152) );
  DFFRX1 \block_r_reg[5][9]  ( .D(n5289), .CK(clk), .RN(n4286), .QN(n7896) );
  DFFRX1 \block_r_reg[3][9]  ( .D(n5033), .CK(clk), .RN(n4286), .QN(n7640) );
  DFFRX1 \block_r_reg[7][111]  ( .D(n5647), .CK(clk), .RN(n4269), .QN(n8254)
         );
  DFFRX1 \block_r_reg[5][111]  ( .D(n5391), .CK(clk), .RN(n4269), .QN(n7998)
         );
  DFFRX1 \block_r_reg[3][111]  ( .D(n5135), .CK(clk), .RN(n4269), .QN(n7742)
         );
  DFFRX1 \block_r_reg[7][110]  ( .D(n5646), .CK(clk), .RN(n4268), .QN(n8253)
         );
  DFFRX1 \block_r_reg[5][110]  ( .D(n5390), .CK(clk), .RN(n4268), .QN(n7997)
         );
  DFFRX1 \block_r_reg[3][110]  ( .D(n5134), .CK(clk), .RN(n4268), .QN(n7741)
         );
  DFFRX1 \block_r_reg[7][109]  ( .D(n5645), .CK(clk), .RN(n4268), .QN(n8252)
         );
  DFFRX1 \block_r_reg[5][109]  ( .D(n5389), .CK(clk), .RN(n4268), .QN(n7996)
         );
  DFFRX1 \block_r_reg[3][109]  ( .D(n5133), .CK(clk), .RN(n4267), .QN(n7740)
         );
  DFFRX1 \block_r_reg[7][108]  ( .D(n5644), .CK(clk), .RN(n4267), .QN(n8251)
         );
  DFFRX1 \block_r_reg[5][108]  ( .D(n5388), .CK(clk), .RN(n4267), .QN(n7995)
         );
  DFFRX1 \block_r_reg[3][108]  ( .D(n5132), .CK(clk), .RN(n4267), .QN(n7739)
         );
  DFFRX1 \block_r_reg[7][107]  ( .D(n5643), .CK(clk), .RN(n4266), .QN(n8250)
         );
  DFFRX1 \block_r_reg[5][107]  ( .D(n5387), .CK(clk), .RN(n4266), .QN(n7994)
         );
  DFFRX1 \block_r_reg[3][107]  ( .D(n5131), .CK(clk), .RN(n4266), .QN(n7738)
         );
  DFFRX1 \block_r_reg[7][106]  ( .D(n5642), .CK(clk), .RN(n4266), .QN(n8249)
         );
  DFFRX1 \block_r_reg[5][106]  ( .D(n5386), .CK(clk), .RN(n4266), .QN(n7993)
         );
  DFFRX1 \block_r_reg[3][106]  ( .D(n5130), .CK(clk), .RN(n4265), .QN(n7737)
         );
  DFFRX1 \block_r_reg[7][105]  ( .D(n5641), .CK(clk), .RN(n4265), .QN(n8248)
         );
  DFFRX1 \block_r_reg[5][105]  ( .D(n5385), .CK(clk), .RN(n4265), .QN(n7992)
         );
  DFFRX1 \block_r_reg[3][105]  ( .D(n5129), .CK(clk), .RN(n4265), .QN(n7736)
         );
  DFFRX1 \block_r_reg[7][79]  ( .D(n5615), .CK(clk), .RN(n4248), .QN(n8222) );
  DFFRX1 \block_r_reg[5][79]  ( .D(n5359), .CK(clk), .RN(n4248), .QN(n7966) );
  DFFRX1 \block_r_reg[3][79]  ( .D(n5103), .CK(clk), .RN(n4247), .QN(n7710) );
  DFFRX1 \block_r_reg[7][78]  ( .D(n5614), .CK(clk), .RN(n4247), .QN(n8221) );
  DFFRX1 \block_r_reg[5][78]  ( .D(n5358), .CK(clk), .RN(n4247), .QN(n7965) );
  DFFRX1 \block_r_reg[3][78]  ( .D(n5102), .CK(clk), .RN(n4247), .QN(n7709) );
  DFFRX1 \block_r_reg[7][77]  ( .D(n5613), .CK(clk), .RN(n4246), .QN(n8220) );
  DFFRX1 \block_r_reg[5][77]  ( .D(n5357), .CK(clk), .RN(n4246), .QN(n7964) );
  DFFRX1 \block_r_reg[3][77]  ( .D(n5101), .CK(clk), .RN(n4246), .QN(n7708) );
  DFFRX1 \block_r_reg[7][76]  ( .D(n5612), .CK(clk), .RN(n4246), .QN(n8219) );
  DFFRX1 \block_r_reg[5][76]  ( .D(n5356), .CK(clk), .RN(n4246), .QN(n7963) );
  DFFRX1 \block_r_reg[3][76]  ( .D(n5100), .CK(clk), .RN(n4245), .QN(n7707) );
  DFFRX1 \block_r_reg[7][75]  ( .D(n5611), .CK(clk), .RN(n4245), .QN(n8218) );
  DFFRX1 \block_r_reg[5][75]  ( .D(n5355), .CK(clk), .RN(n4245), .QN(n7962) );
  DFFRX1 \block_r_reg[3][75]  ( .D(n5099), .CK(clk), .RN(n4245), .QN(n7706) );
  DFFRX1 \block_r_reg[7][74]  ( .D(n5610), .CK(clk), .RN(n4244), .QN(n8217) );
  DFFRX1 \block_r_reg[5][74]  ( .D(n5354), .CK(clk), .RN(n4244), .QN(n7961) );
  DFFRX1 \block_r_reg[3][74]  ( .D(n5098), .CK(clk), .RN(n4244), .QN(n7705) );
  DFFRX1 \block_r_reg[7][73]  ( .D(n5609), .CK(clk), .RN(n4244), .QN(n8216) );
  DFFRX1 \block_r_reg[5][73]  ( .D(n5353), .CK(clk), .RN(n4244), .QN(n7960) );
  DFFRX1 \block_r_reg[3][73]  ( .D(n5097), .CK(clk), .RN(n4243), .QN(n7704) );
  DFFRX1 \block_r_reg[3][72]  ( .D(n5096), .CK(clk), .RN(n4243), .QN(n7703) );
  DFFRX1 \block_r_reg[7][47]  ( .D(n5583), .CK(clk), .RN(n4226), .QN(n8190) );
  DFFRX1 \block_r_reg[5][47]  ( .D(n5327), .CK(clk), .RN(n4226), .QN(n7934) );
  DFFRX1 \block_r_reg[3][47]  ( .D(n5071), .CK(clk), .RN(n4226), .QN(n7678) );
  DFFRX1 \block_r_reg[7][46]  ( .D(n5582), .CK(clk), .RN(n4226), .QN(n8189) );
  DFFRX1 \block_r_reg[5][46]  ( .D(n5326), .CK(clk), .RN(n4226), .QN(n7933) );
  DFFRX1 \block_r_reg[3][46]  ( .D(n5070), .CK(clk), .RN(n4225), .QN(n7677) );
  DFFRX1 \block_r_reg[7][45]  ( .D(n5581), .CK(clk), .RN(n4225), .QN(n8188) );
  DFFRX1 \block_r_reg[5][45]  ( .D(n5325), .CK(clk), .RN(n4225), .QN(n7932) );
  DFFRX1 \block_r_reg[3][45]  ( .D(n5069), .CK(clk), .RN(n4225), .QN(n7676) );
  DFFRX1 \block_r_reg[7][44]  ( .D(n5580), .CK(clk), .RN(n4224), .QN(n8187) );
  DFFRX1 \block_r_reg[5][44]  ( .D(n5324), .CK(clk), .RN(n4224), .QN(n7931) );
  DFFRX1 \block_r_reg[3][44]  ( .D(n5068), .CK(clk), .RN(n4224), .QN(n7675) );
  DFFRX1 \block_r_reg[7][43]  ( .D(n5579), .CK(clk), .RN(n4224), .QN(n8186) );
  DFFRX1 \block_r_reg[5][43]  ( .D(n5323), .CK(clk), .RN(n4224), .QN(n7930) );
  DFFRX1 \block_r_reg[3][43]  ( .D(n5067), .CK(clk), .RN(n4223), .QN(n7674) );
  DFFRX1 \block_r_reg[7][42]  ( .D(n5578), .CK(clk), .RN(n4223), .QN(n8185) );
  DFFRX1 \block_r_reg[5][42]  ( .D(n5322), .CK(clk), .RN(n4223), .QN(n7929) );
  DFFRX1 \block_r_reg[3][42]  ( .D(n5066), .CK(clk), .RN(n4223), .QN(n7673) );
  DFFRX1 \block_r_reg[7][41]  ( .D(n5577), .CK(clk), .RN(n4222), .QN(n8184) );
  DFFRX1 \block_r_reg[5][41]  ( .D(n5321), .CK(clk), .RN(n4222), .QN(n7928) );
  DFFRX1 \block_r_reg[3][41]  ( .D(n5065), .CK(clk), .RN(n4222), .QN(n7672) );
  DFFRX1 \block_r_reg[3][40]  ( .D(n5064), .CK(clk), .RN(n4221), .QN(n7671) );
  DFFRX1 \block_r_reg[0][15]  ( .D(n4655), .CK(clk), .RN(n4290), .QN(n7262) );
  DFFRX1 \block_r_reg[6][15]  ( .D(n5423), .CK(clk), .RN(n4290), .QN(n8030) );
  DFFRX1 \block_r_reg[4][15]  ( .D(n5167), .CK(clk), .RN(n4290), .QN(n7774) );
  DFFRX1 \block_r_reg[2][15]  ( .D(n4911), .CK(clk), .RN(n4290), .QN(n7518) );
  DFFRX1 \block_r_reg[0][14]  ( .D(n4654), .CK(clk), .RN(n4290), .QN(n7261) );
  DFFRX1 \block_r_reg[6][14]  ( .D(n5422), .CK(clk), .RN(n4290), .QN(n8029) );
  DFFRX1 \block_r_reg[4][14]  ( .D(n5166), .CK(clk), .RN(n4289), .QN(n7773) );
  DFFRX1 \block_r_reg[2][14]  ( .D(n4910), .CK(clk), .RN(n4289), .QN(n7517) );
  DFFRX1 \block_r_reg[0][13]  ( .D(n4653), .CK(clk), .RN(n4289), .QN(n7260) );
  DFFRX1 \block_r_reg[6][13]  ( .D(n5421), .CK(clk), .RN(n4289), .QN(n8028) );
  DFFRX1 \block_r_reg[4][13]  ( .D(n5165), .CK(clk), .RN(n4289), .QN(n7772) );
  DFFRX1 \block_r_reg[2][13]  ( .D(n4909), .CK(clk), .RN(n4289), .QN(n7516) );
  DFFRX1 \block_r_reg[0][12]  ( .D(n4652), .CK(clk), .RN(n4288), .QN(n7259) );
  DFFRX1 \block_r_reg[6][12]  ( .D(n5420), .CK(clk), .RN(n4288), .QN(n8027) );
  DFFRX1 \block_r_reg[4][12]  ( .D(n5164), .CK(clk), .RN(n4288), .QN(n7771) );
  DFFRX1 \block_r_reg[2][12]  ( .D(n4908), .CK(clk), .RN(n4288), .QN(n7515) );
  DFFRX1 \block_r_reg[0][11]  ( .D(n4651), .CK(clk), .RN(n4288), .QN(n7258) );
  DFFRX1 \block_r_reg[6][11]  ( .D(n5419), .CK(clk), .RN(n4288), .QN(n8026) );
  DFFRX1 \block_r_reg[4][11]  ( .D(n5163), .CK(clk), .RN(n4287), .QN(n7770) );
  DFFRX1 \block_r_reg[2][11]  ( .D(n4907), .CK(clk), .RN(n4287), .QN(n7514) );
  DFFRX1 \block_r_reg[0][10]  ( .D(n4650), .CK(clk), .RN(n4287), .QN(n7257) );
  DFFRX1 \block_r_reg[6][10]  ( .D(n5418), .CK(clk), .RN(n4287), .QN(n8025) );
  DFFRX1 \block_r_reg[4][10]  ( .D(n5162), .CK(clk), .RN(n4287), .QN(n7769) );
  DFFRX1 \block_r_reg[2][10]  ( .D(n4906), .CK(clk), .RN(n4287), .QN(n7513) );
  DFFRX1 \block_r_reg[0][9]  ( .D(n4649), .CK(clk), .RN(n4286), .QN(n7256) );
  DFFRX1 \block_r_reg[6][9]  ( .D(n5417), .CK(clk), .RN(n4286), .QN(n8024) );
  DFFRX1 \block_r_reg[4][9]  ( .D(n5161), .CK(clk), .RN(n4286), .QN(n7768) );
  DFFRX1 \block_r_reg[2][9]  ( .D(n4905), .CK(clk), .RN(n4286), .QN(n7512) );
  DFFRX1 \block_r_reg[0][111]  ( .D(n4751), .CK(clk), .RN(n4269), .QN(n7358)
         );
  DFFRX1 \block_r_reg[6][111]  ( .D(n5519), .CK(clk), .RN(n4269), .QN(n8126)
         );
  DFFRX1 \block_r_reg[4][111]  ( .D(n5263), .CK(clk), .RN(n4269), .QN(n7870)
         );
  DFFRX1 \block_r_reg[2][111]  ( .D(n5007), .CK(clk), .RN(n4269), .QN(n7614)
         );
  DFFRX1 \block_r_reg[0][110]  ( .D(n4750), .CK(clk), .RN(n4268), .QN(n7357)
         );
  DFFRX1 \block_r_reg[6][110]  ( .D(n5518), .CK(clk), .RN(n4268), .QN(n8125)
         );
  DFFRX1 \block_r_reg[4][110]  ( .D(n5262), .CK(clk), .RN(n4268), .QN(n7869)
         );
  DFFRX1 \block_r_reg[2][110]  ( .D(n5006), .CK(clk), .RN(n4268), .QN(n7613)
         );
  DFFRX1 \block_r_reg[0][109]  ( .D(n4749), .CK(clk), .RN(n4268), .QN(n7356)
         );
  DFFRX1 \block_r_reg[6][109]  ( .D(n5517), .CK(clk), .RN(n4268), .QN(n8124)
         );
  DFFRX1 \block_r_reg[4][109]  ( .D(n5261), .CK(clk), .RN(n4267), .QN(n7868)
         );
  DFFRX1 \block_r_reg[2][109]  ( .D(n5005), .CK(clk), .RN(n4267), .QN(n7612)
         );
  DFFRX1 \block_r_reg[0][108]  ( .D(n4748), .CK(clk), .RN(n4267), .QN(n7355)
         );
  DFFRX1 \block_r_reg[6][108]  ( .D(n5516), .CK(clk), .RN(n4267), .QN(n8123)
         );
  DFFRX1 \block_r_reg[4][108]  ( .D(n5260), .CK(clk), .RN(n4267), .QN(n7867)
         );
  DFFRX1 \block_r_reg[2][108]  ( .D(n5004), .CK(clk), .RN(n4267), .QN(n7611)
         );
  DFFRX1 \block_r_reg[0][107]  ( .D(n4747), .CK(clk), .RN(n4266), .QN(n7354)
         );
  DFFRX1 \block_r_reg[6][107]  ( .D(n5515), .CK(clk), .RN(n4266), .QN(n8122)
         );
  DFFRX1 \block_r_reg[4][107]  ( .D(n5259), .CK(clk), .RN(n4266), .QN(n7866)
         );
  DFFRX1 \block_r_reg[2][107]  ( .D(n5003), .CK(clk), .RN(n4266), .QN(n7610)
         );
  DFFRX1 \block_r_reg[0][106]  ( .D(n4746), .CK(clk), .RN(n4266), .QN(n7353)
         );
  DFFRX1 \block_r_reg[6][106]  ( .D(n5514), .CK(clk), .RN(n4266), .QN(n8121)
         );
  DFFRX1 \block_r_reg[4][106]  ( .D(n5258), .CK(clk), .RN(n4265), .QN(n7865)
         );
  DFFRX1 \block_r_reg[2][106]  ( .D(n5002), .CK(clk), .RN(n4265), .QN(n7609)
         );
  DFFRX1 \block_r_reg[0][105]  ( .D(n4745), .CK(clk), .RN(n4265), .QN(n7352)
         );
  DFFRX1 \block_r_reg[6][105]  ( .D(n5513), .CK(clk), .RN(n4265), .QN(n8120)
         );
  DFFRX1 \block_r_reg[4][105]  ( .D(n5257), .CK(clk), .RN(n4265), .QN(n7864)
         );
  DFFRX1 \block_r_reg[2][105]  ( .D(n5001), .CK(clk), .RN(n4265), .QN(n7608)
         );
  DFFRX1 \block_r_reg[0][79]  ( .D(n4719), .CK(clk), .RN(n4248), .QN(n7326) );
  DFFRX1 \block_r_reg[6][79]  ( .D(n5487), .CK(clk), .RN(n4248), .QN(n8094) );
  DFFRX1 \block_r_reg[4][79]  ( .D(n5231), .CK(clk), .RN(n4247), .QN(n7838) );
  DFFRX1 \block_r_reg[2][79]  ( .D(n4975), .CK(clk), .RN(n4247), .QN(n7582) );
  DFFRX1 \block_r_reg[0][78]  ( .D(n4718), .CK(clk), .RN(n4247), .QN(n7325) );
  DFFRX1 \block_r_reg[6][78]  ( .D(n5486), .CK(clk), .RN(n4247), .QN(n8093) );
  DFFRX1 \block_r_reg[4][78]  ( .D(n5230), .CK(clk), .RN(n4247), .QN(n7837) );
  DFFRX1 \block_r_reg[2][78]  ( .D(n4974), .CK(clk), .RN(n4247), .QN(n7581) );
  DFFRX1 \block_r_reg[0][77]  ( .D(n4717), .CK(clk), .RN(n4246), .QN(n7324) );
  DFFRX1 \block_r_reg[6][77]  ( .D(n5485), .CK(clk), .RN(n4246), .QN(n8092) );
  DFFRX1 \block_r_reg[4][77]  ( .D(n5229), .CK(clk), .RN(n4246), .QN(n7836) );
  DFFRX1 \block_r_reg[2][77]  ( .D(n4973), .CK(clk), .RN(n4246), .QN(n7580) );
  DFFRX1 \block_r_reg[0][76]  ( .D(n4716), .CK(clk), .RN(n4246), .QN(n7323) );
  DFFRX1 \block_r_reg[6][76]  ( .D(n5484), .CK(clk), .RN(n4246), .QN(n8091) );
  DFFRX1 \block_r_reg[4][76]  ( .D(n5228), .CK(clk), .RN(n4245), .QN(n7835) );
  DFFRX1 \block_r_reg[2][76]  ( .D(n4972), .CK(clk), .RN(n4245), .QN(n7579) );
  DFFRX1 \block_r_reg[0][75]  ( .D(n4715), .CK(clk), .RN(n4245), .QN(n7322) );
  DFFRX1 \block_r_reg[6][75]  ( .D(n5483), .CK(clk), .RN(n4245), .QN(n8090) );
  DFFRX1 \block_r_reg[4][75]  ( .D(n5227), .CK(clk), .RN(n4245), .QN(n7834) );
  DFFRX1 \block_r_reg[2][75]  ( .D(n4971), .CK(clk), .RN(n4245), .QN(n7578) );
  DFFRX1 \block_r_reg[0][74]  ( .D(n4714), .CK(clk), .RN(n4244), .QN(n7321) );
  DFFRX1 \block_r_reg[6][74]  ( .D(n5482), .CK(clk), .RN(n4244), .QN(n8089) );
  DFFRX1 \block_r_reg[4][74]  ( .D(n5226), .CK(clk), .RN(n4244), .QN(n7833) );
  DFFRX1 \block_r_reg[2][74]  ( .D(n4970), .CK(clk), .RN(n4244), .QN(n7577) );
  DFFRX1 \block_r_reg[0][73]  ( .D(n4713), .CK(clk), .RN(n4244), .QN(n7320) );
  DFFRX1 \block_r_reg[6][73]  ( .D(n5481), .CK(clk), .RN(n4244), .QN(n8088) );
  DFFRX1 \block_r_reg[4][73]  ( .D(n5225), .CK(clk), .RN(n4243), .QN(n7832) );
  DFFRX1 \block_r_reg[2][73]  ( .D(n4969), .CK(clk), .RN(n4243), .QN(n7576) );
  DFFRX1 \block_r_reg[0][72]  ( .D(n4712), .CK(clk), .RN(n4243), .QN(n7319) );
  DFFRX1 \block_r_reg[2][72]  ( .D(n4968), .CK(clk), .RN(n4243), .QN(n7575) );
  DFFRX1 \block_r_reg[0][47]  ( .D(n4687), .CK(clk), .RN(n4226), .QN(n7294) );
  DFFRX1 \block_r_reg[6][47]  ( .D(n5455), .CK(clk), .RN(n4226), .QN(n8062) );
  DFFRX1 \block_r_reg[4][47]  ( .D(n5199), .CK(clk), .RN(n4226), .QN(n7806) );
  DFFRX1 \block_r_reg[2][47]  ( .D(n4943), .CK(clk), .RN(n4226), .QN(n7550) );
  DFFRX1 \block_r_reg[0][46]  ( .D(n4686), .CK(clk), .RN(n4226), .QN(n7293) );
  DFFRX1 \block_r_reg[6][46]  ( .D(n5454), .CK(clk), .RN(n4226), .QN(n8061) );
  DFFRX1 \block_r_reg[4][46]  ( .D(n5198), .CK(clk), .RN(n4225), .QN(n7805) );
  DFFRX1 \block_r_reg[2][46]  ( .D(n4942), .CK(clk), .RN(n4225), .QN(n7549) );
  DFFRX1 \block_r_reg[0][45]  ( .D(n4685), .CK(clk), .RN(n4225), .QN(n7292) );
  DFFRX1 \block_r_reg[6][45]  ( .D(n5453), .CK(clk), .RN(n4225), .QN(n8060) );
  DFFRX1 \block_r_reg[4][45]  ( .D(n5197), .CK(clk), .RN(n4225), .QN(n7804) );
  DFFRX1 \block_r_reg[2][45]  ( .D(n4941), .CK(clk), .RN(n4225), .QN(n7548) );
  DFFRX1 \block_r_reg[0][44]  ( .D(n4684), .CK(clk), .RN(n4224), .QN(n7291) );
  DFFRX1 \block_r_reg[6][44]  ( .D(n5452), .CK(clk), .RN(n4224), .QN(n8059) );
  DFFRX1 \block_r_reg[4][44]  ( .D(n5196), .CK(clk), .RN(n4224), .QN(n7803) );
  DFFRX1 \block_r_reg[2][44]  ( .D(n4940), .CK(clk), .RN(n4224), .QN(n7547) );
  DFFRX1 \block_r_reg[0][43]  ( .D(n4683), .CK(clk), .RN(n4224), .QN(n7290) );
  DFFRX1 \block_r_reg[6][43]  ( .D(n5451), .CK(clk), .RN(n4224), .QN(n8058) );
  DFFRX1 \block_r_reg[4][43]  ( .D(n5195), .CK(clk), .RN(n4223), .QN(n7802) );
  DFFRX1 \block_r_reg[2][43]  ( .D(n4939), .CK(clk), .RN(n4223), .QN(n7546) );
  DFFRX1 \block_r_reg[0][42]  ( .D(n4682), .CK(clk), .RN(n4223), .QN(n7289) );
  DFFRX1 \block_r_reg[6][42]  ( .D(n5450), .CK(clk), .RN(n4223), .QN(n8057) );
  DFFRX1 \block_r_reg[4][42]  ( .D(n5194), .CK(clk), .RN(n4223), .QN(n7801) );
  DFFRX1 \block_r_reg[2][42]  ( .D(n4938), .CK(clk), .RN(n4223), .QN(n7545) );
  DFFRX1 \block_r_reg[0][41]  ( .D(n4681), .CK(clk), .RN(n4222), .QN(n7288) );
  DFFRX1 \block_r_reg[6][41]  ( .D(n5449), .CK(clk), .RN(n4222), .QN(n8056) );
  DFFRX1 \block_r_reg[4][41]  ( .D(n5193), .CK(clk), .RN(n4222), .QN(n7800) );
  DFFRX1 \block_r_reg[2][41]  ( .D(n4937), .CK(clk), .RN(n4222), .QN(n7544) );
  DFFRX1 \block_r_reg[0][40]  ( .D(n4680), .CK(clk), .RN(n4222), .QN(n7287) );
  DFFRX1 \block_r_reg[6][40]  ( .D(n5448), .CK(clk), .RN(n4222), .QN(n8055) );
  DFFRX1 \block_r_reg[2][40]  ( .D(n4936), .CK(clk), .RN(n4221), .QN(n7543) );
  DFFRX1 \tag_r_reg[1][24]  ( .D(n4615), .CK(clk), .RN(n4308), .Q(n1302), .QN(
        n7096) );
  DFFRX1 \tag_r_reg[1][23]  ( .D(n4614), .CK(clk), .RN(n4308), .QN(n7095) );
  DFFRX1 \tag_r_reg[1][22]  ( .D(n4613), .CK(clk), .RN(n4308), .QN(n7094) );
  DFFRX1 \tag_r_reg[1][21]  ( .D(n4612), .CK(clk), .RN(n4308), .QN(n7093) );
  DFFRX1 \tag_r_reg[1][20]  ( .D(n4611), .CK(clk), .RN(n4308), .QN(n7092) );
  DFFRX1 \tag_r_reg[1][19]  ( .D(n4610), .CK(clk), .RN(n4308), .QN(n7091) );
  DFFRX1 \tag_r_reg[1][11]  ( .D(n4602), .CK(clk), .RN(n4307), .QN(n7083) );
  DFFRX1 \tag_r_reg[1][10]  ( .D(n4601), .CK(clk), .RN(n4307), .QN(n7082) );
  DFFRX1 \tag_r_reg[1][9]  ( .D(n4600), .CK(clk), .RN(n4307), .QN(n7081) );
  DFFRX1 \tag_r_reg[1][8]  ( .D(n4599), .CK(clk), .RN(n4307), .QN(n7080) );
  DFFRX1 \tag_r_reg[1][7]  ( .D(n4598), .CK(clk), .RN(n4307), .QN(n7079) );
  DFFRX1 \tag_r_reg[1][5]  ( .D(n4596), .CK(clk), .RN(n4307), .QN(n7077) );
  DFFRX1 \tag_r_reg[3][24]  ( .D(n4565), .CK(clk), .RN(n4304), .Q(n1300), .QN(
        n7146) );
  DFFRX1 \tag_r_reg[3][23]  ( .D(n4564), .CK(clk), .RN(n4304), .QN(n7145) );
  DFFRX1 \tag_r_reg[3][22]  ( .D(n4563), .CK(clk), .RN(n4304), .QN(n7144) );
  DFFRX1 \tag_r_reg[3][21]  ( .D(n4562), .CK(clk), .RN(n4304), .QN(n7143) );
  DFFRX1 \tag_r_reg[3][20]  ( .D(n4561), .CK(clk), .RN(n4304), .QN(n7142) );
  DFFRX1 \tag_r_reg[3][19]  ( .D(n4560), .CK(clk), .RN(n4304), .QN(n7141) );
  DFFRX1 \tag_r_reg[3][9]  ( .D(n4550), .CK(clk), .RN(n4303), .QN(n7131) );
  DFFRX1 \tag_r_reg[3][8]  ( .D(n4549), .CK(clk), .RN(n4303), .QN(n7130) );
  DFFRX1 \tag_r_reg[3][7]  ( .D(n4548), .CK(clk), .RN(n4303), .QN(n7129) );
  DFFRX1 \tag_r_reg[5][24]  ( .D(n4515), .CK(clk), .RN(n4300), .Q(n1303), .QN(
        n7196) );
  DFFRX1 \tag_r_reg[5][23]  ( .D(n4514), .CK(clk), .RN(n4300), .QN(n7195) );
  DFFRX1 \tag_r_reg[5][22]  ( .D(n4513), .CK(clk), .RN(n4300), .QN(n7194) );
  DFFRX1 \tag_r_reg[5][21]  ( .D(n4512), .CK(clk), .RN(n4300), .QN(n7193) );
  DFFRX1 \tag_r_reg[5][20]  ( .D(n4511), .CK(clk), .RN(n4300), .QN(n7192) );
  DFFRX1 \tag_r_reg[5][19]  ( .D(n4510), .CK(clk), .RN(n4300), .QN(n7191) );
  DFFRX1 \tag_r_reg[5][11]  ( .D(n4502), .CK(clk), .RN(n4299), .QN(n7183) );
  DFFRX1 \tag_r_reg[5][10]  ( .D(n4501), .CK(clk), .RN(n4299), .QN(n7182) );
  DFFRX1 \tag_r_reg[5][9]  ( .D(n4500), .CK(clk), .RN(n4299), .QN(n7181) );
  DFFRX1 \tag_r_reg[5][8]  ( .D(n4499), .CK(clk), .RN(n4299), .QN(n7180) );
  DFFRX1 \tag_r_reg[5][7]  ( .D(n4498), .CK(clk), .RN(n4299), .QN(n7179) );
  DFFRX1 \tag_r_reg[5][5]  ( .D(n4496), .CK(clk), .RN(n4298), .QN(n7177) );
  DFFRX1 \tag_r_reg[7][24]  ( .D(n4465), .CK(clk), .RN(n4296), .Q(n1298), .QN(
        n7246) );
  DFFRX1 \tag_r_reg[7][23]  ( .D(n4464), .CK(clk), .RN(n4296), .QN(n7245) );
  DFFRX1 \tag_r_reg[7][22]  ( .D(n4463), .CK(clk), .RN(n4296), .QN(n7244) );
  DFFRX1 \tag_r_reg[7][21]  ( .D(n4462), .CK(clk), .RN(n4296), .QN(n7243) );
  DFFRX1 \tag_r_reg[7][20]  ( .D(n4461), .CK(clk), .RN(n4296), .QN(n7242) );
  DFFRX1 \tag_r_reg[7][19]  ( .D(n4460), .CK(clk), .RN(n4295), .QN(n7241) );
  DFFRX1 \tag_r_reg[7][9]  ( .D(n4450), .CK(clk), .RN(n4295), .QN(n7231) );
  DFFRX1 \tag_r_reg[7][8]  ( .D(n4449), .CK(clk), .RN(n4295), .QN(n7230) );
  DFFRX1 \tag_r_reg[7][7]  ( .D(n4448), .CK(clk), .RN(n4294), .QN(n7229) );
  DFFRX1 \tag_r_reg[2][24]  ( .D(n4590), .CK(clk), .RN(n4306), .Q(n1301), .QN(
        n7121) );
  DFFRX1 \tag_r_reg[2][23]  ( .D(n4589), .CK(clk), .RN(n4306), .QN(n7120) );
  DFFRX1 \tag_r_reg[2][22]  ( .D(n4588), .CK(clk), .RN(n4306), .QN(n7119) );
  DFFRX1 \tag_r_reg[2][21]  ( .D(n4587), .CK(clk), .RN(n4306), .QN(n7118) );
  DFFRX1 \tag_r_reg[2][20]  ( .D(n4586), .CK(clk), .RN(n4306), .QN(n7117) );
  DFFRX1 \tag_r_reg[2][19]  ( .D(n4585), .CK(clk), .RN(n4306), .QN(n7116) );
  DFFRX1 \tag_r_reg[2][10]  ( .D(n4576), .CK(clk), .RN(n4305), .QN(n7107) );
  DFFRX1 \tag_r_reg[2][9]  ( .D(n4575), .CK(clk), .RN(n4305), .QN(n7106) );
  DFFRX1 \tag_r_reg[2][8]  ( .D(n4574), .CK(clk), .RN(n4305), .QN(n7105) );
  DFFRX1 \tag_r_reg[2][7]  ( .D(n4573), .CK(clk), .RN(n4305), .QN(n7104) );
  DFFRX1 \tag_r_reg[4][24]  ( .D(n4540), .CK(clk), .RN(n4302), .Q(n1304), .QN(
        n7171) );
  DFFRX1 \tag_r_reg[4][23]  ( .D(n4539), .CK(clk), .RN(n4302), .QN(n7170) );
  DFFRX1 \tag_r_reg[4][22]  ( .D(n4538), .CK(clk), .RN(n4302), .QN(n7169) );
  DFFRX1 \tag_r_reg[4][21]  ( .D(n4537), .CK(clk), .RN(n4302), .QN(n7168) );
  DFFRX1 \tag_r_reg[4][20]  ( .D(n4536), .CK(clk), .RN(n4302), .QN(n7167) );
  DFFRX1 \tag_r_reg[4][19]  ( .D(n4535), .CK(clk), .RN(n4302), .QN(n7166) );
  DFFRX1 \tag_r_reg[4][11]  ( .D(n4527), .CK(clk), .RN(n4301), .QN(n7158) );
  DFFRX1 \tag_r_reg[4][10]  ( .D(n4526), .CK(clk), .RN(n4301), .QN(n7157) );
  DFFRX1 \tag_r_reg[4][9]  ( .D(n4525), .CK(clk), .RN(n4301), .QN(n7156) );
  DFFRX1 \tag_r_reg[4][8]  ( .D(n4524), .CK(clk), .RN(n4301), .QN(n7155) );
  DFFRX1 \tag_r_reg[4][7]  ( .D(n4523), .CK(clk), .RN(n4301), .QN(n7154) );
  DFFRX1 \tag_r_reg[4][5]  ( .D(n4521), .CK(clk), .RN(n4301), .QN(n7152) );
  DFFRX1 \tag_r_reg[6][24]  ( .D(n4490), .CK(clk), .RN(n4298), .Q(n1299), .QN(
        n7221) );
  DFFRX1 \tag_r_reg[6][23]  ( .D(n4489), .CK(clk), .RN(n4298), .QN(n7220) );
  DFFRX1 \tag_r_reg[6][22]  ( .D(n4488), .CK(clk), .RN(n4298), .QN(n7219) );
  DFFRX1 \tag_r_reg[6][21]  ( .D(n4487), .CK(clk), .RN(n4298), .QN(n7218) );
  DFFRX1 \tag_r_reg[6][20]  ( .D(n4486), .CK(clk), .RN(n4298), .QN(n7217) );
  DFFRX1 \tag_r_reg[6][19]  ( .D(n4485), .CK(clk), .RN(n4298), .QN(n7216) );
  DFFRX1 \tag_r_reg[6][11]  ( .D(n4477), .CK(clk), .RN(n4297), .QN(n7208) );
  DFFRX1 \tag_r_reg[6][10]  ( .D(n4476), .CK(clk), .RN(n4297), .QN(n7207) );
  DFFRX1 \tag_r_reg[6][9]  ( .D(n4475), .CK(clk), .RN(n4297), .QN(n7206) );
  DFFRX1 \tag_r_reg[6][8]  ( .D(n4474), .CK(clk), .RN(n4297), .QN(n7205) );
  DFFRX1 \tag_r_reg[6][7]  ( .D(n4473), .CK(clk), .RN(n4297), .QN(n7204) );
  DFFRX1 \tag_r_reg[6][5]  ( .D(n4471), .CK(clk), .RN(n4296), .QN(n7202) );
  DFFRX1 \tag_r_reg[0][24]  ( .D(n4639), .CK(clk), .RN(n4294), .Q(n1297), .QN(
        n7071) );
  DFFRX1 \tag_r_reg[0][23]  ( .D(n4638), .CK(clk), .RN(n4294), .QN(n7070) );
  DFFRX1 \tag_r_reg[0][22]  ( .D(n4637), .CK(clk), .RN(n4294), .QN(n7069) );
  DFFRX1 \tag_r_reg[0][21]  ( .D(n4636), .CK(clk), .RN(n4294), .QN(n7068) );
  DFFRX1 \tag_r_reg[0][20]  ( .D(n4635), .CK(clk), .RN(n4293), .QN(n7067) );
  DFFRX1 \tag_r_reg[0][19]  ( .D(n4634), .CK(clk), .RN(n4293), .QN(n7066) );
  DFFRX1 \tag_r_reg[0][16]  ( .D(n4631), .CK(clk), .RN(n4293), .QN(n7063) );
  DFFRX1 \tag_r_reg[0][10]  ( .D(n4625), .CK(clk), .RN(n4293), .QN(n7057) );
  DFFRX1 \tag_r_reg[0][9]  ( .D(n4624), .CK(clk), .RN(n4293), .QN(n7056) );
  DFFRX1 \tag_r_reg[0][8]  ( .D(n4623), .CK(clk), .RN(n4292), .QN(n7055) );
  DFFRX1 \tag_r_reg[0][7]  ( .D(n4622), .CK(clk), .RN(n4292), .QN(n7054) );
  DFFRX1 \tag_r_reg[0][5]  ( .D(n4620), .CK(clk), .RN(n4292), .QN(n7052) );
  DFFRX1 \block_r_reg[1][8]  ( .D(n4776), .CK(clk), .RN(n4285), .QN(n7383) );
  DFFRX1 \block_r_reg[1][7]  ( .D(n4775), .CK(clk), .RN(n4285), .QN(n7382) );
  DFFRX1 \block_r_reg[1][6]  ( .D(n4774), .CK(clk), .RN(n4284), .QN(n7381) );
  DFFRX1 \block_r_reg[5][5]  ( .D(n5285), .CK(clk), .RN(n4284), .QN(n7892) );
  DFFRX1 \block_r_reg[1][5]  ( .D(n4773), .CK(clk), .RN(n4283), .QN(n7380) );
  DFFRX1 \block_r_reg[5][4]  ( .D(n5284), .CK(clk), .RN(n4283), .QN(n7891) );
  DFFRX1 \block_r_reg[1][4]  ( .D(n4772), .CK(clk), .RN(n4283), .QN(n7379) );
  DFFRX1 \block_r_reg[5][3]  ( .D(n5283), .CK(clk), .RN(n4282), .QN(n7890) );
  DFFRX1 \block_r_reg[1][3]  ( .D(n4771), .CK(clk), .RN(n4282), .QN(n7378) );
  DFFRX1 \block_r_reg[5][2]  ( .D(n5282), .CK(clk), .RN(n4282), .QN(n7889) );
  DFFRX1 \block_r_reg[1][2]  ( .D(n4770), .CK(clk), .RN(n4281), .QN(n7377) );
  DFFRX1 \block_r_reg[1][1]  ( .D(n4769), .CK(clk), .RN(n4281), .QN(n7376) );
  DFFRX1 \block_r_reg[5][104]  ( .D(n5384), .CK(clk), .RN(n4264), .QN(n7991)
         );
  DFFRX1 \block_r_reg[1][104]  ( .D(n4872), .CK(clk), .RN(n4264), .QN(n7479)
         );
  DFFRX1 \block_r_reg[5][103]  ( .D(n5383), .CK(clk), .RN(n4264), .QN(n7990)
         );
  DFFRX1 \block_r_reg[1][103]  ( .D(n4871), .CK(clk), .RN(n4263), .QN(n7478)
         );
  DFFRX1 \block_r_reg[5][102]  ( .D(n5382), .CK(clk), .RN(n4263), .QN(n7989)
         );
  DFFRX1 \block_r_reg[1][102]  ( .D(n4870), .CK(clk), .RN(n4263), .QN(n7477)
         );
  DFFRX1 \block_r_reg[5][101]  ( .D(n5381), .CK(clk), .RN(n4262), .QN(n7988)
         );
  DFFRX1 \block_r_reg[1][101]  ( .D(n4869), .CK(clk), .RN(n4262), .QN(n7476)
         );
  DFFRX1 \block_r_reg[5][100]  ( .D(n5380), .CK(clk), .RN(n4262), .QN(n7987)
         );
  DFFRX1 \block_r_reg[1][100]  ( .D(n4868), .CK(clk), .RN(n4261), .QN(n7475)
         );
  DFFRX1 \block_r_reg[5][99]  ( .D(n5379), .CK(clk), .RN(n4261), .QN(n7986) );
  DFFRX1 \block_r_reg[1][99]  ( .D(n4867), .CK(clk), .RN(n4261), .QN(n7474) );
  DFFRX1 \block_r_reg[5][98]  ( .D(n5378), .CK(clk), .RN(n4260), .QN(n7985) );
  DFFRX1 \block_r_reg[1][98]  ( .D(n4866), .CK(clk), .RN(n4260), .QN(n7473) );
  DFFRX1 \block_r_reg[1][97]  ( .D(n4865), .CK(clk), .RN(n4259), .QN(n7472) );
  DFFRX1 \block_r_reg[1][71]  ( .D(n4839), .CK(clk), .RN(n4242), .QN(n7446) );
  DFFRX1 \block_r_reg[1][70]  ( .D(n4838), .CK(clk), .RN(n4241), .QN(n7445) );
  DFFRX1 \block_r_reg[1][69]  ( .D(n4837), .CK(clk), .RN(n4241), .QN(n7444) );
  DFFRX1 \block_r_reg[1][68]  ( .D(n4836), .CK(clk), .RN(n4240), .QN(n7443) );
  DFFRX1 \block_r_reg[1][67]  ( .D(n4835), .CK(clk), .RN(n4239), .QN(n7442) );
  DFFRX1 \block_r_reg[1][66]  ( .D(n4834), .CK(clk), .RN(n4239), .QN(n7441) );
  DFFRX1 \block_r_reg[1][65]  ( .D(n4833), .CK(clk), .RN(n4238), .QN(n7440) );
  DFFRX1 \block_r_reg[1][64]  ( .D(n4832), .CK(clk), .RN(n4237), .QN(n7439) );
  DFFRX1 \block_r_reg[1][39]  ( .D(n4807), .CK(clk), .RN(n4221), .QN(n7414) );
  DFFRX1 \block_r_reg[1][38]  ( .D(n4806), .CK(clk), .RN(n4220), .QN(n7413) );
  DFFRX1 \block_r_reg[1][37]  ( .D(n4805), .CK(clk), .RN(n4219), .QN(n7412) );
  DFFRX1 \block_r_reg[1][36]  ( .D(n4804), .CK(clk), .RN(n4219), .QN(n7411) );
  DFFRX1 \block_r_reg[1][35]  ( .D(n4803), .CK(clk), .RN(n4218), .QN(n7410) );
  DFFRX1 \block_r_reg[1][34]  ( .D(n4802), .CK(clk), .RN(n4217), .QN(n7409) );
  DFFRX1 \block_r_reg[1][33]  ( .D(n4801), .CK(clk), .RN(n4217), .QN(n7408) );
  DFFRX1 \block_r_reg[1][32]  ( .D(n4800), .CK(clk), .RN(n4216), .QN(n7407) );
  DFFRX1 \block_r_reg[7][8]  ( .D(n5544), .CK(clk), .RN(n4286), .QN(n8151) );
  DFFRX1 \block_r_reg[5][8]  ( .D(n5288), .CK(clk), .RN(n4286), .QN(n7895) );
  DFFRX1 \block_r_reg[3][8]  ( .D(n5032), .CK(clk), .RN(n4285), .QN(n7639) );
  DFFRX1 \block_r_reg[7][7]  ( .D(n5543), .CK(clk), .RN(n4285), .QN(n8150) );
  DFFRX1 \block_r_reg[5][7]  ( .D(n5287), .CK(clk), .RN(n4285), .QN(n7894) );
  DFFRX1 \block_r_reg[3][7]  ( .D(n5031), .CK(clk), .RN(n4285), .QN(n7638) );
  DFFRX1 \block_r_reg[7][6]  ( .D(n5542), .CK(clk), .RN(n4284), .QN(n8149) );
  DFFRX1 \block_r_reg[5][6]  ( .D(n5286), .CK(clk), .RN(n4284), .QN(n7893) );
  DFFRX1 \block_r_reg[3][6]  ( .D(n5030), .CK(clk), .RN(n4284), .QN(n7637) );
  DFFRX1 \block_r_reg[7][5]  ( .D(n5541), .CK(clk), .RN(n4284), .QN(n8148) );
  DFFRX1 \block_r_reg[3][5]  ( .D(n5029), .CK(clk), .RN(n4283), .QN(n7636) );
  DFFRX1 \block_r_reg[7][4]  ( .D(n5540), .CK(clk), .RN(n4283), .QN(n8147) );
  DFFRX1 \block_r_reg[3][4]  ( .D(n5028), .CK(clk), .RN(n4283), .QN(n7635) );
  DFFRX1 \block_r_reg[7][3]  ( .D(n5539), .CK(clk), .RN(n4282), .QN(n8146) );
  DFFRX1 \block_r_reg[3][3]  ( .D(n5027), .CK(clk), .RN(n4282), .QN(n7634) );
  DFFRX1 \block_r_reg[7][2]  ( .D(n5538), .CK(clk), .RN(n4282), .QN(n8145) );
  DFFRX1 \block_r_reg[3][2]  ( .D(n5026), .CK(clk), .RN(n4281), .QN(n7633) );
  DFFRX1 \block_r_reg[7][1]  ( .D(n5537), .CK(clk), .RN(n4281), .QN(n8144) );
  DFFRX1 \block_r_reg[3][1]  ( .D(n5025), .CK(clk), .RN(n4281), .QN(n7632) );
  DFFRX1 \block_r_reg[7][104]  ( .D(n5640), .CK(clk), .RN(n4264), .QN(n8247)
         );
  DFFRX1 \block_r_reg[3][104]  ( .D(n5128), .CK(clk), .RN(n4264), .QN(n7735)
         );
  DFFRX1 \block_r_reg[7][103]  ( .D(n5639), .CK(clk), .RN(n4264), .QN(n8246)
         );
  DFFRX1 \block_r_reg[3][103]  ( .D(n5127), .CK(clk), .RN(n4263), .QN(n7734)
         );
  DFFRX1 \block_r_reg[7][102]  ( .D(n5638), .CK(clk), .RN(n4263), .QN(n8245)
         );
  DFFRX1 \block_r_reg[3][102]  ( .D(n5126), .CK(clk), .RN(n4263), .QN(n7733)
         );
  DFFRX1 \block_r_reg[7][101]  ( .D(n5637), .CK(clk), .RN(n4262), .QN(n8244)
         );
  DFFRX1 \block_r_reg[3][101]  ( .D(n5125), .CK(clk), .RN(n4262), .QN(n7732)
         );
  DFFRX1 \block_r_reg[7][100]  ( .D(n5636), .CK(clk), .RN(n4262), .QN(n8243)
         );
  DFFRX1 \block_r_reg[3][100]  ( .D(n5124), .CK(clk), .RN(n4261), .QN(n7731)
         );
  DFFRX1 \block_r_reg[7][99]  ( .D(n5635), .CK(clk), .RN(n4261), .QN(n8242) );
  DFFRX1 \block_r_reg[3][99]  ( .D(n5123), .CK(clk), .RN(n4261), .QN(n7730) );
  DFFRX1 \block_r_reg[7][98]  ( .D(n5634), .CK(clk), .RN(n4260), .QN(n8241) );
  DFFRX1 \block_r_reg[3][98]  ( .D(n5122), .CK(clk), .RN(n4260), .QN(n7729) );
  DFFRX1 \block_r_reg[7][97]  ( .D(n5633), .CK(clk), .RN(n4260), .QN(n8240) );
  DFFRX1 \block_r_reg[3][97]  ( .D(n5121), .CK(clk), .RN(n4259), .QN(n7728) );
  DFFRX1 \block_r_reg[7][72]  ( .D(n5608), .CK(clk), .RN(n4243), .QN(n8215) );
  DFFRX1 \block_r_reg[5][72]  ( .D(n5352), .CK(clk), .RN(n4243), .QN(n7959) );
  DFFRX1 \block_r_reg[7][71]  ( .D(n5607), .CK(clk), .RN(n4242), .QN(n8214) );
  DFFRX1 \block_r_reg[5][71]  ( .D(n5351), .CK(clk), .RN(n4242), .QN(n7958) );
  DFFRX1 \block_r_reg[3][71]  ( .D(n5095), .CK(clk), .RN(n4242), .QN(n7702) );
  DFFRX1 \block_r_reg[7][70]  ( .D(n5606), .CK(clk), .RN(n4242), .QN(n8213) );
  DFFRX1 \block_r_reg[5][70]  ( .D(n5350), .CK(clk), .RN(n4242), .QN(n7957) );
  DFFRX1 \block_r_reg[3][70]  ( .D(n5094), .CK(clk), .RN(n4241), .QN(n7701) );
  DFFRX1 \block_r_reg[7][69]  ( .D(n5605), .CK(clk), .RN(n4241), .QN(n8212) );
  DFFRX1 \block_r_reg[5][69]  ( .D(n5349), .CK(clk), .RN(n4241), .QN(n7956) );
  DFFRX1 \block_r_reg[3][69]  ( .D(n5093), .CK(clk), .RN(n4241), .QN(n7700) );
  DFFRX1 \block_r_reg[7][68]  ( .D(n5604), .CK(clk), .RN(n4240), .QN(n8211) );
  DFFRX1 \block_r_reg[5][68]  ( .D(n5348), .CK(clk), .RN(n4240), .QN(n7955) );
  DFFRX1 \block_r_reg[3][68]  ( .D(n5092), .CK(clk), .RN(n4240), .QN(n7699) );
  DFFRX1 \block_r_reg[7][67]  ( .D(n5603), .CK(clk), .RN(n4240), .QN(n8210) );
  DFFRX1 \block_r_reg[5][67]  ( .D(n5347), .CK(clk), .RN(n4240), .QN(n7954) );
  DFFRX1 \block_r_reg[3][67]  ( .D(n5091), .CK(clk), .RN(n4239), .QN(n7698) );
  DFFRX1 \block_r_reg[7][66]  ( .D(n5602), .CK(clk), .RN(n4239), .QN(n8209) );
  DFFRX1 \block_r_reg[5][66]  ( .D(n5346), .CK(clk), .RN(n4239), .QN(n7953) );
  DFFRX1 \block_r_reg[3][66]  ( .D(n5090), .CK(clk), .RN(n4239), .QN(n7697) );
  DFFRX1 \block_r_reg[7][65]  ( .D(n5601), .CK(clk), .RN(n4238), .QN(n8208) );
  DFFRX1 \block_r_reg[5][65]  ( .D(n5345), .CK(clk), .RN(n4238), .QN(n7952) );
  DFFRX1 \block_r_reg[3][65]  ( .D(n5089), .CK(clk), .RN(n4238), .QN(n7696) );
  DFFRX1 \block_r_reg[7][64]  ( .D(n5600), .CK(clk), .RN(n4238), .QN(n8207) );
  DFFRX1 \block_r_reg[5][64]  ( .D(n5344), .CK(clk), .RN(n4238), .QN(n7951) );
  DFFRX1 \block_r_reg[3][64]  ( .D(n5088), .CK(clk), .RN(n4237), .QN(n7695) );
  DFFRX1 \block_r_reg[7][40]  ( .D(n5576), .CK(clk), .RN(n4222), .QN(n8183) );
  DFFRX1 \block_r_reg[5][40]  ( .D(n5320), .CK(clk), .RN(n4222), .QN(n7927) );
  DFFRX1 \block_r_reg[7][39]  ( .D(n5575), .CK(clk), .RN(n4221), .QN(n8182) );
  DFFRX1 \block_r_reg[5][39]  ( .D(n5319), .CK(clk), .RN(n4221), .QN(n7926) );
  DFFRX1 \block_r_reg[3][39]  ( .D(n5063), .CK(clk), .RN(n4221), .QN(n7670) );
  DFFRX1 \block_r_reg[7][38]  ( .D(n5574), .CK(clk), .RN(n4220), .QN(n8181) );
  DFFRX1 \block_r_reg[5][38]  ( .D(n5318), .CK(clk), .RN(n4220), .QN(n7925) );
  DFFRX1 \block_r_reg[3][38]  ( .D(n5062), .CK(clk), .RN(n4220), .QN(n7669) );
  DFFRX1 \block_r_reg[7][37]  ( .D(n5573), .CK(clk), .RN(n4220), .QN(n8180) );
  DFFRX1 \block_r_reg[5][37]  ( .D(n5317), .CK(clk), .RN(n4220), .QN(n7924) );
  DFFRX1 \block_r_reg[3][37]  ( .D(n5061), .CK(clk), .RN(n4219), .QN(n7668) );
  DFFRX1 \block_r_reg[7][36]  ( .D(n5572), .CK(clk), .RN(n4219), .QN(n8179) );
  DFFRX1 \block_r_reg[5][36]  ( .D(n5316), .CK(clk), .RN(n4219), .QN(n7923) );
  DFFRX1 \block_r_reg[3][36]  ( .D(n5060), .CK(clk), .RN(n4219), .QN(n7667) );
  DFFRX1 \block_r_reg[7][35]  ( .D(n5571), .CK(clk), .RN(n4218), .QN(n8178) );
  DFFRX1 \block_r_reg[5][35]  ( .D(n5315), .CK(clk), .RN(n4218), .QN(n7922) );
  DFFRX1 \block_r_reg[3][35]  ( .D(n5059), .CK(clk), .RN(n4218), .QN(n7666) );
  DFFRX1 \block_r_reg[7][34]  ( .D(n5570), .CK(clk), .RN(n4218), .QN(n8177) );
  DFFRX1 \block_r_reg[5][34]  ( .D(n5314), .CK(clk), .RN(n4218), .QN(n7921) );
  DFFRX1 \block_r_reg[4][34]  ( .D(n5186), .CK(clk), .RN(n4217), .QN(n7793) );
  DFFRX1 \block_r_reg[3][34]  ( .D(n5058), .CK(clk), .RN(n4217), .QN(n7665) );
  DFFRX1 \block_r_reg[7][33]  ( .D(n5569), .CK(clk), .RN(n4217), .QN(n8176) );
  DFFRX1 \block_r_reg[5][33]  ( .D(n5313), .CK(clk), .RN(n4217), .QN(n7920) );
  DFFRX1 \block_r_reg[4][33]  ( .D(n5185), .CK(clk), .RN(n4217), .QN(n7792) );
  DFFRX1 \block_r_reg[3][33]  ( .D(n5057), .CK(clk), .RN(n4217), .QN(n7664) );
  DFFRX1 \block_r_reg[7][32]  ( .D(n5568), .CK(clk), .RN(n4216), .QN(n8175) );
  DFFRX1 \block_r_reg[5][32]  ( .D(n5312), .CK(clk), .RN(n4216), .QN(n7919) );
  DFFRX1 \block_r_reg[4][32]  ( .D(n5184), .CK(clk), .RN(n4216), .QN(n7791) );
  DFFRX1 \block_r_reg[3][32]  ( .D(n5056), .CK(clk), .RN(n4216), .QN(n7663) );
  DFFRX1 \block_r_reg[0][8]  ( .D(n4648), .CK(clk), .RN(n4286), .QN(n7255) );
  DFFRX1 \block_r_reg[6][8]  ( .D(n5416), .CK(clk), .RN(n4286), .QN(n8023) );
  DFFRX1 \block_r_reg[4][8]  ( .D(n5160), .CK(clk), .RN(n4285), .QN(n7767) );
  DFFRX1 \block_r_reg[2][8]  ( .D(n4904), .CK(clk), .RN(n4285), .QN(n7511) );
  DFFRX1 \block_r_reg[0][7]  ( .D(n4647), .CK(clk), .RN(n4285), .QN(n7254) );
  DFFRX1 \block_r_reg[6][7]  ( .D(n5415), .CK(clk), .RN(n4285), .QN(n8022) );
  DFFRX1 \block_r_reg[4][7]  ( .D(n5159), .CK(clk), .RN(n4285), .QN(n7766) );
  DFFRX1 \block_r_reg[2][7]  ( .D(n4903), .CK(clk), .RN(n4285), .QN(n7510) );
  DFFRX1 \block_r_reg[0][6]  ( .D(n4646), .CK(clk), .RN(n4284), .QN(n7253) );
  DFFRX1 \block_r_reg[6][6]  ( .D(n5414), .CK(clk), .RN(n4284), .QN(n8021) );
  DFFRX1 \block_r_reg[4][6]  ( .D(n5158), .CK(clk), .RN(n4284), .QN(n7765) );
  DFFRX1 \block_r_reg[2][6]  ( .D(n4902), .CK(clk), .RN(n4284), .QN(n7509) );
  DFFRX1 \block_r_reg[0][5]  ( .D(n4645), .CK(clk), .RN(n4284), .QN(n7252) );
  DFFRX1 \block_r_reg[6][5]  ( .D(n5413), .CK(clk), .RN(n4284), .QN(n8020) );
  DFFRX1 \block_r_reg[4][5]  ( .D(n5157), .CK(clk), .RN(n4283), .QN(n7764) );
  DFFRX1 \block_r_reg[2][5]  ( .D(n4901), .CK(clk), .RN(n4283), .QN(n7508) );
  DFFRX1 \block_r_reg[0][4]  ( .D(n4644), .CK(clk), .RN(n4283), .QN(n7251) );
  DFFRX1 \block_r_reg[6][4]  ( .D(n5412), .CK(clk), .RN(n4283), .QN(n8019) );
  DFFRX1 \block_r_reg[4][4]  ( .D(n5156), .CK(clk), .RN(n4283), .QN(n7763) );
  DFFRX1 \block_r_reg[2][4]  ( .D(n4900), .CK(clk), .RN(n4283), .QN(n7507) );
  DFFRX1 \block_r_reg[0][3]  ( .D(n4643), .CK(clk), .RN(n4282), .QN(n7250) );
  DFFRX1 \block_r_reg[6][3]  ( .D(n5411), .CK(clk), .RN(n4282), .QN(n8018) );
  DFFRX1 \block_r_reg[4][3]  ( .D(n5155), .CK(clk), .RN(n4282), .QN(n7762) );
  DFFRX1 \block_r_reg[2][3]  ( .D(n4899), .CK(clk), .RN(n4282), .QN(n7506) );
  DFFRX1 \block_r_reg[0][2]  ( .D(n4642), .CK(clk), .RN(n4282), .QN(n7249) );
  DFFRX1 \block_r_reg[6][2]  ( .D(n5410), .CK(clk), .RN(n4282), .QN(n8017) );
  DFFRX1 \block_r_reg[4][2]  ( .D(n5154), .CK(clk), .RN(n4281), .QN(n7761) );
  DFFRX1 \block_r_reg[2][2]  ( .D(n4898), .CK(clk), .RN(n4281), .QN(n7505) );
  DFFRX1 \block_r_reg[0][1]  ( .D(n4641), .CK(clk), .RN(n4281), .QN(n7248) );
  DFFRX1 \block_r_reg[6][1]  ( .D(n5409), .CK(clk), .RN(n4281), .QN(n8016) );
  DFFRX1 \block_r_reg[4][1]  ( .D(n5153), .CK(clk), .RN(n4281), .QN(n7760) );
  DFFRX1 \block_r_reg[2][1]  ( .D(n4897), .CK(clk), .RN(n4281), .QN(n7504) );
  DFFRX1 \block_r_reg[2][0]  ( .D(n4896), .CK(clk), .RN(n4280), .QN(n7503) );
  DFFRX1 \block_r_reg[0][104]  ( .D(n4744), .CK(clk), .RN(n4264), .QN(n7351)
         );
  DFFRX1 \block_r_reg[6][104]  ( .D(n5512), .CK(clk), .RN(n4264), .QN(n8119)
         );
  DFFRX1 \block_r_reg[4][104]  ( .D(n5256), .CK(clk), .RN(n4264), .QN(n7863)
         );
  DFFRX1 \block_r_reg[2][104]  ( .D(n5000), .CK(clk), .RN(n4264), .QN(n7607)
         );
  DFFRX1 \block_r_reg[0][103]  ( .D(n4743), .CK(clk), .RN(n4264), .QN(n7350)
         );
  DFFRX1 \block_r_reg[6][103]  ( .D(n5511), .CK(clk), .RN(n4264), .QN(n8118)
         );
  DFFRX1 \block_r_reg[4][103]  ( .D(n5255), .CK(clk), .RN(n4263), .QN(n7862)
         );
  DFFRX1 \block_r_reg[2][103]  ( .D(n4999), .CK(clk), .RN(n4263), .QN(n7606)
         );
  DFFRX1 \block_r_reg[0][102]  ( .D(n4742), .CK(clk), .RN(n4263), .QN(n7349)
         );
  DFFRX1 \block_r_reg[6][102]  ( .D(n5510), .CK(clk), .RN(n4263), .QN(n8117)
         );
  DFFRX1 \block_r_reg[4][102]  ( .D(n5254), .CK(clk), .RN(n4263), .QN(n7861)
         );
  DFFRX1 \block_r_reg[2][102]  ( .D(n4998), .CK(clk), .RN(n4263), .QN(n7605)
         );
  DFFRX1 \block_r_reg[0][101]  ( .D(n4741), .CK(clk), .RN(n4262), .QN(n7348)
         );
  DFFRX1 \block_r_reg[6][101]  ( .D(n5509), .CK(clk), .RN(n4262), .QN(n8116)
         );
  DFFRX1 \block_r_reg[4][101]  ( .D(n5253), .CK(clk), .RN(n4262), .QN(n7860)
         );
  DFFRX1 \block_r_reg[2][101]  ( .D(n4997), .CK(clk), .RN(n4262), .QN(n7604)
         );
  DFFRX1 \block_r_reg[0][100]  ( .D(n4740), .CK(clk), .RN(n4262), .QN(n7347)
         );
  DFFRX1 \block_r_reg[6][100]  ( .D(n5508), .CK(clk), .RN(n4262), .QN(n8115)
         );
  DFFRX1 \block_r_reg[4][100]  ( .D(n5252), .CK(clk), .RN(n4261), .QN(n7859)
         );
  DFFRX1 \block_r_reg[2][100]  ( .D(n4996), .CK(clk), .RN(n4261), .QN(n7603)
         );
  DFFRX1 \block_r_reg[0][99]  ( .D(n4739), .CK(clk), .RN(n4261), .QN(n7346) );
  DFFRX1 \block_r_reg[6][99]  ( .D(n5507), .CK(clk), .RN(n4261), .QN(n8114) );
  DFFRX1 \block_r_reg[4][99]  ( .D(n5251), .CK(clk), .RN(n4261), .QN(n7858) );
  DFFRX1 \block_r_reg[2][99]  ( .D(n4995), .CK(clk), .RN(n4261), .QN(n7602) );
  DFFRX1 \block_r_reg[0][98]  ( .D(n4738), .CK(clk), .RN(n4260), .QN(n7345) );
  DFFRX1 \block_r_reg[6][98]  ( .D(n5506), .CK(clk), .RN(n4260), .QN(n8113) );
  DFFRX1 \block_r_reg[4][98]  ( .D(n5250), .CK(clk), .RN(n4260), .QN(n7857) );
  DFFRX1 \block_r_reg[2][98]  ( .D(n4994), .CK(clk), .RN(n4260), .QN(n7601) );
  DFFRX1 \block_r_reg[0][97]  ( .D(n4737), .CK(clk), .RN(n4260), .QN(n7344) );
  DFFRX1 \block_r_reg[6][97]  ( .D(n5505), .CK(clk), .RN(n4260), .QN(n8112) );
  DFFRX1 \block_r_reg[2][97]  ( .D(n4993), .CK(clk), .RN(n4259), .QN(n7600) );
  DFFRX1 \block_r_reg[6][72]  ( .D(n5480), .CK(clk), .RN(n4243), .QN(n8087) );
  DFFRX1 \block_r_reg[4][72]  ( .D(n5224), .CK(clk), .RN(n4243), .QN(n7831) );
  DFFRX1 \block_r_reg[0][71]  ( .D(n4711), .CK(clk), .RN(n4242), .QN(n7318) );
  DFFRX1 \block_r_reg[6][71]  ( .D(n5479), .CK(clk), .RN(n4242), .QN(n8086) );
  DFFRX1 \block_r_reg[4][71]  ( .D(n5223), .CK(clk), .RN(n4242), .QN(n7830) );
  DFFRX1 \block_r_reg[2][71]  ( .D(n4967), .CK(clk), .RN(n4242), .QN(n7574) );
  DFFRX1 \block_r_reg[0][70]  ( .D(n4710), .CK(clk), .RN(n4242), .QN(n7317) );
  DFFRX1 \block_r_reg[6][70]  ( .D(n5478), .CK(clk), .RN(n4242), .QN(n8085) );
  DFFRX1 \block_r_reg[4][70]  ( .D(n5222), .CK(clk), .RN(n4241), .QN(n7829) );
  DFFRX1 \block_r_reg[2][70]  ( .D(n4966), .CK(clk), .RN(n4241), .QN(n7573) );
  DFFRX1 \block_r_reg[0][69]  ( .D(n4709), .CK(clk), .RN(n4241), .QN(n7316) );
  DFFRX1 \block_r_reg[6][69]  ( .D(n5477), .CK(clk), .RN(n4241), .QN(n8084) );
  DFFRX1 \block_r_reg[4][69]  ( .D(n5221), .CK(clk), .RN(n4241), .QN(n7828) );
  DFFRX1 \block_r_reg[2][69]  ( .D(n4965), .CK(clk), .RN(n4241), .QN(n7572) );
  DFFRX1 \block_r_reg[0][68]  ( .D(n4708), .CK(clk), .RN(n4240), .QN(n7315) );
  DFFRX1 \block_r_reg[6][68]  ( .D(n5476), .CK(clk), .RN(n4240), .QN(n8083) );
  DFFRX1 \block_r_reg[4][68]  ( .D(n5220), .CK(clk), .RN(n4240), .QN(n7827) );
  DFFRX1 \block_r_reg[2][68]  ( .D(n4964), .CK(clk), .RN(n4240), .QN(n7571) );
  DFFRX1 \block_r_reg[0][67]  ( .D(n4707), .CK(clk), .RN(n4240), .QN(n7314) );
  DFFRX1 \block_r_reg[6][67]  ( .D(n5475), .CK(clk), .RN(n4240), .QN(n8082) );
  DFFRX1 \block_r_reg[4][67]  ( .D(n5219), .CK(clk), .RN(n4239), .QN(n7826) );
  DFFRX1 \block_r_reg[2][67]  ( .D(n4963), .CK(clk), .RN(n4239), .QN(n7570) );
  DFFRX1 \block_r_reg[0][66]  ( .D(n4706), .CK(clk), .RN(n4239), .QN(n7313) );
  DFFRX1 \block_r_reg[6][66]  ( .D(n5474), .CK(clk), .RN(n4239), .QN(n8081) );
  DFFRX1 \block_r_reg[4][66]  ( .D(n5218), .CK(clk), .RN(n4239), .QN(n7825) );
  DFFRX1 \block_r_reg[2][66]  ( .D(n4962), .CK(clk), .RN(n4239), .QN(n7569) );
  DFFRX1 \block_r_reg[0][65]  ( .D(n4705), .CK(clk), .RN(n4238), .QN(n7312) );
  DFFRX1 \block_r_reg[6][65]  ( .D(n5473), .CK(clk), .RN(n4238), .QN(n8080) );
  DFFRX1 \block_r_reg[4][65]  ( .D(n5217), .CK(clk), .RN(n4238), .QN(n7824) );
  DFFRX1 \block_r_reg[2][65]  ( .D(n4961), .CK(clk), .RN(n4238), .QN(n7568) );
  DFFRX1 \block_r_reg[0][64]  ( .D(n4704), .CK(clk), .RN(n4238), .QN(n7311) );
  DFFRX1 \block_r_reg[6][64]  ( .D(n5472), .CK(clk), .RN(n4238), .QN(n8079) );
  DFFRX1 \block_r_reg[4][64]  ( .D(n5216), .CK(clk), .RN(n4237), .QN(n7823) );
  DFFRX1 \block_r_reg[2][64]  ( .D(n4960), .CK(clk), .RN(n4237), .QN(n7567) );
  DFFRX1 \block_r_reg[4][40]  ( .D(n5192), .CK(clk), .RN(n4221), .QN(n7799) );
  DFFRX1 \block_r_reg[0][39]  ( .D(n4679), .CK(clk), .RN(n4221), .QN(n7286) );
  DFFRX1 \block_r_reg[6][39]  ( .D(n5447), .CK(clk), .RN(n4221), .QN(n8054) );
  DFFRX1 \block_r_reg[4][39]  ( .D(n5191), .CK(clk), .RN(n4221), .QN(n7798) );
  DFFRX1 \block_r_reg[2][39]  ( .D(n4935), .CK(clk), .RN(n4221), .QN(n7542) );
  DFFRX1 \block_r_reg[0][38]  ( .D(n4678), .CK(clk), .RN(n4220), .QN(n7285) );
  DFFRX1 \block_r_reg[6][38]  ( .D(n5446), .CK(clk), .RN(n4220), .QN(n8053) );
  DFFRX1 \block_r_reg[4][38]  ( .D(n5190), .CK(clk), .RN(n4220), .QN(n7797) );
  DFFRX1 \block_r_reg[2][38]  ( .D(n4934), .CK(clk), .RN(n4220), .QN(n7541) );
  DFFRX1 \block_r_reg[0][37]  ( .D(n4677), .CK(clk), .RN(n4220), .QN(n7284) );
  DFFRX1 \block_r_reg[6][37]  ( .D(n5445), .CK(clk), .RN(n4220), .QN(n8052) );
  DFFRX1 \block_r_reg[4][37]  ( .D(n5189), .CK(clk), .RN(n4219), .QN(n7796) );
  DFFRX1 \block_r_reg[2][37]  ( .D(n4933), .CK(clk), .RN(n4219), .QN(n7540) );
  DFFRX1 \block_r_reg[0][36]  ( .D(n4676), .CK(clk), .RN(n4219), .QN(n7283) );
  DFFRX1 \block_r_reg[6][36]  ( .D(n5444), .CK(clk), .RN(n4219), .QN(n8051) );
  DFFRX1 \block_r_reg[4][36]  ( .D(n5188), .CK(clk), .RN(n4219), .QN(n7795) );
  DFFRX1 \block_r_reg[2][36]  ( .D(n4932), .CK(clk), .RN(n4219), .QN(n7539) );
  DFFRX1 \block_r_reg[0][35]  ( .D(n4675), .CK(clk), .RN(n4218), .QN(n7282) );
  DFFRX1 \block_r_reg[6][35]  ( .D(n5443), .CK(clk), .RN(n4218), .QN(n8050) );
  DFFRX1 \block_r_reg[4][35]  ( .D(n5187), .CK(clk), .RN(n4218), .QN(n7794) );
  DFFRX1 \block_r_reg[2][35]  ( .D(n4931), .CK(clk), .RN(n4218), .QN(n7538) );
  DFFRX1 \block_r_reg[0][34]  ( .D(n4674), .CK(clk), .RN(n4218), .QN(n7281) );
  DFFRX1 \block_r_reg[6][34]  ( .D(n5442), .CK(clk), .RN(n4218), .QN(n8049) );
  DFFRX1 \block_r_reg[2][34]  ( .D(n4930), .CK(clk), .RN(n4217), .QN(n7537) );
  DFFRX1 \block_r_reg[0][33]  ( .D(n4673), .CK(clk), .RN(n4217), .QN(n7280) );
  DFFRX1 \block_r_reg[6][33]  ( .D(n5441), .CK(clk), .RN(n4217), .QN(n8048) );
  DFFRX1 \block_r_reg[2][33]  ( .D(n4929), .CK(clk), .RN(n4217), .QN(n7536) );
  DFFRX1 \block_r_reg[0][32]  ( .D(n4672), .CK(clk), .RN(n4216), .QN(n7279) );
  DFFRX1 \block_r_reg[6][32]  ( .D(n5440), .CK(clk), .RN(n4216), .QN(n8047) );
  DFFRX1 \block_r_reg[2][32]  ( .D(n4928), .CK(clk), .RN(n4216), .QN(n7535) );
  DFFRX1 \block_r_reg[5][1]  ( .D(n5281), .CK(clk), .RN(n4281), .QN(n7888) );
  DFFRX1 \block_r_reg[5][0]  ( .D(n5280), .CK(clk), .RN(n4280), .QN(n7887) );
  DFFRX1 \block_r_reg[1][0]  ( .D(n4768), .CK(clk), .RN(n4280), .QN(n7375) );
  DFFRX1 \block_r_reg[5][97]  ( .D(n5377), .CK(clk), .RN(n4260), .QN(n7984) );
  DFFRX1 \block_r_reg[5][96]  ( .D(n5376), .CK(clk), .RN(n4259), .QN(n7983) );
  DFFRX1 \block_r_reg[1][96]  ( .D(n4864), .CK(clk), .RN(n4259), .QN(n7471) );
  DFFRX1 \block_r_reg[7][0]  ( .D(n5536), .CK(clk), .RN(n4280), .QN(n8143) );
  DFFRX1 \block_r_reg[3][0]  ( .D(n5024), .CK(clk), .RN(n4280), .QN(n7631) );
  DFFRX1 \block_r_reg[7][96]  ( .D(n5632), .CK(clk), .RN(n4259), .QN(n8239) );
  DFFRX1 \block_r_reg[3][96]  ( .D(n5120), .CK(clk), .RN(n4259), .QN(n7727) );
  DFFRX1 \block_r_reg[0][0]  ( .D(n4640), .CK(clk), .RN(n4280), .QN(n7247) );
  DFFRX1 \block_r_reg[6][0]  ( .D(n5408), .CK(clk), .RN(n4280), .QN(n8015) );
  DFFRX1 \block_r_reg[4][0]  ( .D(n5152), .CK(clk), .RN(n4280), .QN(n7759) );
  DFFRX1 \block_r_reg[4][97]  ( .D(n5249), .CK(clk), .RN(n4259), .QN(n7856) );
  DFFRX1 \block_r_reg[0][96]  ( .D(n4736), .CK(clk), .RN(n4259), .QN(n7343) );
  DFFRX1 \block_r_reg[6][96]  ( .D(n5504), .CK(clk), .RN(n4259), .QN(n8111) );
  DFFRX1 \block_r_reg[4][96]  ( .D(n5248), .CK(clk), .RN(n4259), .QN(n7855) );
  DFFRX1 \block_r_reg[2][96]  ( .D(n4992), .CK(clk), .RN(n4259), .QN(n7599) );
  DFFRX1 \state_r_reg[0]  ( .D(n4424), .CK(clk), .RN(n4310), .Q(\state_r[0] ), 
        .QN(n8271) );
  DFFRX1 \state_r_reg[1]  ( .D(n4423), .CK(clk), .RN(n4310), .Q(n8289), .QN(
        n8272) );
  OAI221X1 U3 ( .A0(n6980), .A1(n4204), .B0(n6979), .B1(n4200), .C0(n6978), 
        .Y(proc_rdata[27]) );
  OAI221X1 U4 ( .A0(n6985), .A1(n4205), .B0(n6984), .B1(n4200), .C0(n6983), 
        .Y(proc_rdata[28]) );
  NAND2X1 U5 ( .A(n1333), .B(n6830), .Y(n1) );
  NAND2X1 U6 ( .A(n1333), .B(n4132), .Y(n2) );
  CLKBUFX2 U7 ( .A(n6712), .Y(n4053) );
  NAND2X1 U8 ( .A(n1333), .B(n4142), .Y(n3) );
  NAND2X1 U9 ( .A(n1333), .B(n4152), .Y(n4) );
  CLKBUFX2 U10 ( .A(n6713), .Y(n4060) );
  NAND2X1 U11 ( .A(n1333), .B(n6856), .Y(n5) );
  NAND2X1 U12 ( .A(n1333), .B(n6854), .Y(n6) );
  NAND2X1 U13 ( .A(n1333), .B(n6858), .Y(n7) );
  CLKBUFX2 U14 ( .A(n6710), .Y(n4024) );
  NAND2X1 U15 ( .A(n1333), .B(n4122), .Y(n8) );
  NAND2X1 U16 ( .A(n8289), .B(n8271), .Y(n9) );
  OA22X1 U17 ( .A0(n4003), .A1(n4402), .B0(n5788), .B1(n4004), .Y(n10) );
  OA22X1 U18 ( .A0(n4003), .A1(n4412), .B0(n5713), .B1(n4004), .Y(n11) );
  OA22X1 U19 ( .A0(n4003), .A1(n4413), .B0(n5718), .B1(n4004), .Y(n12) );
  OA22X1 U20 ( .A0(n4003), .A1(n4414), .B0(n5723), .B1(n4005), .Y(n13) );
  OA22X1 U21 ( .A0(n4003), .A1(n4415), .B0(n5728), .B1(n4005), .Y(n14) );
  OA22X1 U22 ( .A0(n4003), .A1(n4416), .B0(n5733), .B1(n4005), .Y(n15) );
  OA22X1 U23 ( .A0(n4003), .A1(n4419), .B0(n5748), .B1(n4004), .Y(n16) );
  OA22X1 U24 ( .A0(n4003), .A1(n4420), .B0(n5753), .B1(n4005), .Y(n17) );
  OA22X1 U25 ( .A0(n4003), .A1(n4417), .B0(n5738), .B1(n4005), .Y(n18) );
  OA22X1 U26 ( .A0(n4003), .A1(n4418), .B0(n5743), .B1(n4005), .Y(n19) );
  INVX12 U27 ( .A(n6882), .Y(mem_wdata[0]) );
  NOR4X2 U28 ( .A(n5792), .B(n5791), .C(n5790), .D(n5789), .Y(n6882) );
  INVX12 U29 ( .A(n7011), .Y(mem_wdata[100]) );
  NOR4X2 U30 ( .A(n5796), .B(n5795), .C(n5794), .D(n5793), .Y(n7011) );
  INVX12 U31 ( .A(n7016), .Y(mem_wdata[101]) );
  NOR4X2 U32 ( .A(n5800), .B(n5799), .C(n5798), .D(n5797), .Y(n7016) );
  INVX12 U33 ( .A(n7021), .Y(mem_wdata[102]) );
  NOR4X2 U34 ( .A(n5804), .B(n5803), .C(n5802), .D(n5801), .Y(n7021) );
  INVX12 U35 ( .A(n7026), .Y(mem_wdata[103]) );
  NOR4X2 U36 ( .A(n5808), .B(n5807), .C(n5806), .D(n5805), .Y(n7026) );
  INVX12 U37 ( .A(n7031), .Y(mem_wdata[104]) );
  NOR4X2 U38 ( .A(n5812), .B(n5811), .C(n5810), .D(n5809), .Y(n7031) );
  INVX12 U39 ( .A(n7037), .Y(mem_wdata[105]) );
  NOR4X2 U40 ( .A(n5816), .B(n5815), .C(n5814), .D(n5813), .Y(n7037) );
  INVX12 U41 ( .A(n6886), .Y(mem_wdata[106]) );
  NOR4X2 U42 ( .A(n5820), .B(n5819), .C(n5818), .D(n5817), .Y(n6886) );
  INVX12 U43 ( .A(n6891), .Y(mem_wdata[107]) );
  NOR4X2 U44 ( .A(n5824), .B(n5823), .C(n5822), .D(n5821), .Y(n6891) );
  INVX12 U45 ( .A(n6896), .Y(mem_wdata[108]) );
  NOR4X2 U46 ( .A(n5828), .B(n5827), .C(n5826), .D(n5825), .Y(n6896) );
  INVX12 U47 ( .A(n6901), .Y(mem_wdata[109]) );
  NOR4X2 U48 ( .A(n5832), .B(n5831), .C(n5830), .D(n5829), .Y(n6901) );
  INVX12 U49 ( .A(n6887), .Y(mem_wdata[10]) );
  NOR4X2 U50 ( .A(n5836), .B(n5835), .C(n5834), .D(n5833), .Y(n6887) );
  INVX12 U51 ( .A(n6906), .Y(mem_wdata[110]) );
  NOR4X2 U52 ( .A(n5840), .B(n5839), .C(n5838), .D(n5837), .Y(n6906) );
  INVX12 U53 ( .A(n6911), .Y(mem_wdata[111]) );
  NOR4X2 U54 ( .A(n5844), .B(n5843), .C(n5842), .D(n5841), .Y(n6911) );
  INVX12 U55 ( .A(n6916), .Y(mem_wdata[112]) );
  NOR4X2 U56 ( .A(n5848), .B(n5847), .C(n5846), .D(n5845), .Y(n6916) );
  INVX12 U57 ( .A(n6921), .Y(mem_wdata[113]) );
  NOR4X2 U58 ( .A(n5852), .B(n5851), .C(n5850), .D(n5849), .Y(n6921) );
  INVX12 U59 ( .A(n6926), .Y(mem_wdata[114]) );
  NOR4X2 U60 ( .A(n5856), .B(n5855), .C(n5854), .D(n5853), .Y(n6926) );
  INVX12 U61 ( .A(n6931), .Y(mem_wdata[115]) );
  NOR4X2 U62 ( .A(n5860), .B(n5859), .C(n5858), .D(n5857), .Y(n6931) );
  INVX12 U63 ( .A(n6941), .Y(mem_wdata[116]) );
  NOR4X2 U64 ( .A(n5864), .B(n5863), .C(n5862), .D(n5861), .Y(n6941) );
  INVX12 U65 ( .A(n6946), .Y(mem_wdata[117]) );
  NOR4X2 U66 ( .A(n5868), .B(n5867), .C(n5866), .D(n5865), .Y(n6946) );
  INVX12 U67 ( .A(n6951), .Y(mem_wdata[118]) );
  NOR4X2 U68 ( .A(n5872), .B(n5871), .C(n5870), .D(n5869), .Y(n6951) );
  INVX12 U69 ( .A(n6956), .Y(mem_wdata[119]) );
  NOR4X2 U70 ( .A(n5876), .B(n5875), .C(n5874), .D(n5873), .Y(n6956) );
  INVX12 U71 ( .A(n6892), .Y(mem_wdata[11]) );
  NOR4X2 U72 ( .A(n5880), .B(n5879), .C(n5878), .D(n5877), .Y(n6892) );
  INVX12 U73 ( .A(n6961), .Y(mem_wdata[120]) );
  NOR4X2 U74 ( .A(n5884), .B(n5883), .C(n5882), .D(n5881), .Y(n6961) );
  INVX12 U75 ( .A(n6966), .Y(mem_wdata[121]) );
  NOR4X2 U76 ( .A(n5888), .B(n5887), .C(n5886), .D(n5885), .Y(n6966) );
  INVX12 U77 ( .A(n6971), .Y(mem_wdata[122]) );
  NOR4X2 U78 ( .A(n5892), .B(n5891), .C(n5890), .D(n5889), .Y(n6971) );
  INVX12 U79 ( .A(n6976), .Y(mem_wdata[123]) );
  NOR4X2 U80 ( .A(n5896), .B(n5895), .C(n5894), .D(n5893), .Y(n6976) );
  INVX12 U81 ( .A(n6981), .Y(mem_wdata[124]) );
  NOR4X2 U82 ( .A(n5900), .B(n5899), .C(n5898), .D(n5897), .Y(n6981) );
  INVX12 U83 ( .A(n6986), .Y(mem_wdata[125]) );
  NOR4X2 U84 ( .A(n5904), .B(n5903), .C(n5902), .D(n5901), .Y(n6986) );
  INVX12 U85 ( .A(n6996), .Y(mem_wdata[126]) );
  NOR4X2 U86 ( .A(n5908), .B(n5907), .C(n5906), .D(n5905), .Y(n6996) );
  INVX12 U87 ( .A(n7001), .Y(mem_wdata[127]) );
  NOR4X2 U88 ( .A(n5912), .B(n5911), .C(n5910), .D(n5909), .Y(n7001) );
  INVX12 U89 ( .A(n6897), .Y(mem_wdata[12]) );
  NOR4X2 U90 ( .A(n5916), .B(n5915), .C(n5914), .D(n5913), .Y(n6897) );
  INVX12 U91 ( .A(n6902), .Y(mem_wdata[13]) );
  NOR4X2 U92 ( .A(n5920), .B(n5919), .C(n5918), .D(n5917), .Y(n6902) );
  INVX12 U93 ( .A(n6907), .Y(mem_wdata[14]) );
  NOR4X2 U94 ( .A(n5924), .B(n5923), .C(n5922), .D(n5921), .Y(n6907) );
  INVX12 U95 ( .A(n6912), .Y(mem_wdata[15]) );
  NOR4X2 U96 ( .A(n5928), .B(n5927), .C(n5926), .D(n5925), .Y(n6912) );
  INVX12 U97 ( .A(n6917), .Y(mem_wdata[16]) );
  NOR4X2 U98 ( .A(n5932), .B(n5931), .C(n5930), .D(n5929), .Y(n6917) );
  INVX12 U99 ( .A(n6922), .Y(mem_wdata[17]) );
  NOR4X2 U100 ( .A(n5936), .B(n5935), .C(n5934), .D(n5933), .Y(n6922) );
  INVX12 U101 ( .A(n6927), .Y(mem_wdata[18]) );
  NOR4X2 U102 ( .A(n5940), .B(n5939), .C(n5938), .D(n5937), .Y(n6927) );
  INVX12 U103 ( .A(n6932), .Y(mem_wdata[19]) );
  NOR4X2 U104 ( .A(n5944), .B(n5943), .C(n5942), .D(n5941), .Y(n6932) );
  INVX12 U105 ( .A(n6937), .Y(mem_wdata[1]) );
  NOR4X2 U106 ( .A(n5948), .B(n5947), .C(n5946), .D(n5945), .Y(n6937) );
  INVX12 U107 ( .A(n6942), .Y(mem_wdata[20]) );
  NOR4X2 U108 ( .A(n5952), .B(n5951), .C(n5950), .D(n5949), .Y(n6942) );
  INVX12 U109 ( .A(n6947), .Y(mem_wdata[21]) );
  NOR4X2 U110 ( .A(n5956), .B(n5955), .C(n5954), .D(n5953), .Y(n6947) );
  INVX12 U111 ( .A(n6952), .Y(mem_wdata[22]) );
  NOR4X2 U112 ( .A(n5960), .B(n5959), .C(n5958), .D(n5957), .Y(n6952) );
  INVX12 U113 ( .A(n6957), .Y(mem_wdata[23]) );
  NOR4X2 U114 ( .A(n5964), .B(n5963), .C(n5962), .D(n5961), .Y(n6957) );
  INVX12 U115 ( .A(n6962), .Y(mem_wdata[24]) );
  NOR4X2 U116 ( .A(n5968), .B(n5967), .C(n5966), .D(n5965), .Y(n6962) );
  INVX12 U117 ( .A(n6967), .Y(mem_wdata[25]) );
  NOR4X2 U118 ( .A(n5972), .B(n5971), .C(n5970), .D(n5969), .Y(n6967) );
  INVX12 U119 ( .A(n6972), .Y(mem_wdata[26]) );
  NOR4X2 U120 ( .A(n5976), .B(n5975), .C(n5974), .D(n5973), .Y(n6972) );
  INVX12 U121 ( .A(n6977), .Y(mem_wdata[27]) );
  NOR4X2 U122 ( .A(n5980), .B(n5979), .C(n5978), .D(n5977), .Y(n6977) );
  INVX12 U123 ( .A(n6982), .Y(mem_wdata[28]) );
  NOR4X2 U124 ( .A(n5984), .B(n5983), .C(n5982), .D(n5981), .Y(n6982) );
  INVX12 U125 ( .A(n6987), .Y(mem_wdata[29]) );
  NOR4X2 U126 ( .A(n5988), .B(n5987), .C(n5986), .D(n5985), .Y(n6987) );
  INVX12 U127 ( .A(n6992), .Y(mem_wdata[2]) );
  NOR4X2 U128 ( .A(n5992), .B(n5991), .C(n5990), .D(n5989), .Y(n6992) );
  INVX12 U129 ( .A(n6997), .Y(mem_wdata[30]) );
  NOR4X2 U130 ( .A(n5996), .B(n5995), .C(n5994), .D(n5993), .Y(n6997) );
  INVX12 U131 ( .A(n7002), .Y(mem_wdata[31]) );
  NOR4X2 U132 ( .A(n6000), .B(n5999), .C(n5998), .D(n5997), .Y(n7002) );
  INVX12 U133 ( .A(n6884), .Y(mem_wdata[32]) );
  NOR4X2 U134 ( .A(n6004), .B(n6003), .C(n6002), .D(n6001), .Y(n6884) );
  INVX12 U135 ( .A(n6939), .Y(mem_wdata[33]) );
  NOR4X2 U136 ( .A(n6008), .B(n6007), .C(n6006), .D(n6005), .Y(n6939) );
  INVX12 U137 ( .A(n6994), .Y(mem_wdata[34]) );
  NOR4X2 U138 ( .A(n6012), .B(n6011), .C(n6010), .D(n6009), .Y(n6994) );
  INVX12 U139 ( .A(n7009), .Y(mem_wdata[35]) );
  NOR4X2 U140 ( .A(n6016), .B(n6015), .C(n6014), .D(n6013), .Y(n7009) );
  INVX12 U141 ( .A(n7014), .Y(mem_wdata[36]) );
  NOR4X2 U142 ( .A(n6020), .B(n6019), .C(n6018), .D(n6017), .Y(n7014) );
  INVX12 U143 ( .A(n7019), .Y(mem_wdata[37]) );
  NOR4X2 U144 ( .A(n6024), .B(n6023), .C(n6022), .D(n6021), .Y(n7019) );
  INVX12 U145 ( .A(n7024), .Y(mem_wdata[38]) );
  NOR4X2 U146 ( .A(n6028), .B(n6027), .C(n6026), .D(n6025), .Y(n7024) );
  INVX12 U147 ( .A(n7029), .Y(mem_wdata[39]) );
  NOR4X2 U148 ( .A(n6032), .B(n6031), .C(n6030), .D(n6029), .Y(n7029) );
  INVX12 U149 ( .A(n7007), .Y(mem_wdata[3]) );
  NOR4X2 U150 ( .A(n6036), .B(n6035), .C(n6034), .D(n6033), .Y(n7007) );
  INVX12 U151 ( .A(n7034), .Y(mem_wdata[40]) );
  NOR4X2 U152 ( .A(n6040), .B(n6039), .C(n6038), .D(n6037), .Y(n7034) );
  INVX12 U153 ( .A(n7042), .Y(mem_wdata[41]) );
  NOR4X2 U154 ( .A(n6044), .B(n6043), .C(n6042), .D(n6041), .Y(n7042) );
  INVX12 U155 ( .A(n6889), .Y(mem_wdata[42]) );
  NOR4X2 U156 ( .A(n6048), .B(n6047), .C(n6046), .D(n6045), .Y(n6889) );
  INVX12 U157 ( .A(n6894), .Y(mem_wdata[43]) );
  NOR4X2 U158 ( .A(n6052), .B(n6051), .C(n6050), .D(n6049), .Y(n6894) );
  INVX12 U159 ( .A(n6899), .Y(mem_wdata[44]) );
  NOR4X2 U160 ( .A(n6056), .B(n6055), .C(n6054), .D(n6053), .Y(n6899) );
  INVX12 U161 ( .A(n6904), .Y(mem_wdata[45]) );
  NOR4X2 U162 ( .A(n6060), .B(n6059), .C(n6058), .D(n6057), .Y(n6904) );
  INVX12 U163 ( .A(n6909), .Y(mem_wdata[46]) );
  NOR4X2 U164 ( .A(n6064), .B(n6063), .C(n6062), .D(n6061), .Y(n6909) );
  INVX12 U165 ( .A(n6914), .Y(mem_wdata[47]) );
  NOR4X2 U166 ( .A(n6068), .B(n6067), .C(n6066), .D(n6065), .Y(n6914) );
  INVX12 U167 ( .A(n6919), .Y(mem_wdata[48]) );
  NOR4X2 U168 ( .A(n6072), .B(n6071), .C(n6070), .D(n6069), .Y(n6919) );
  INVX12 U169 ( .A(n6924), .Y(mem_wdata[49]) );
  NOR4X2 U170 ( .A(n6076), .B(n6075), .C(n6074), .D(n6073), .Y(n6924) );
  INVX12 U171 ( .A(n7012), .Y(mem_wdata[4]) );
  NOR4X2 U172 ( .A(n6080), .B(n6079), .C(n6078), .D(n6077), .Y(n7012) );
  INVX12 U173 ( .A(n6929), .Y(mem_wdata[50]) );
  NOR4X2 U174 ( .A(n6084), .B(n6083), .C(n6082), .D(n6081), .Y(n6929) );
  INVX12 U175 ( .A(n6934), .Y(mem_wdata[51]) );
  NOR4X2 U176 ( .A(n6088), .B(n6087), .C(n6086), .D(n6085), .Y(n6934) );
  INVX12 U177 ( .A(n6944), .Y(mem_wdata[52]) );
  NOR4X2 U178 ( .A(n6092), .B(n6091), .C(n6090), .D(n6089), .Y(n6944) );
  INVX12 U179 ( .A(n6949), .Y(mem_wdata[53]) );
  NOR4X2 U180 ( .A(n6096), .B(n6095), .C(n6094), .D(n6093), .Y(n6949) );
  INVX12 U181 ( .A(n6954), .Y(mem_wdata[54]) );
  NOR4X2 U182 ( .A(n6100), .B(n6099), .C(n6098), .D(n6097), .Y(n6954) );
  INVX12 U183 ( .A(n6959), .Y(mem_wdata[55]) );
  NOR4X2 U184 ( .A(n6104), .B(n6103), .C(n6102), .D(n6101), .Y(n6959) );
  INVX12 U185 ( .A(n6964), .Y(mem_wdata[56]) );
  NOR4X2 U186 ( .A(n6108), .B(n6107), .C(n6106), .D(n6105), .Y(n6964) );
  INVX12 U187 ( .A(n6969), .Y(mem_wdata[57]) );
  NOR4X2 U188 ( .A(n6112), .B(n6111), .C(n6110), .D(n6109), .Y(n6969) );
  INVX12 U189 ( .A(n6974), .Y(mem_wdata[58]) );
  NOR4X2 U190 ( .A(n6116), .B(n6115), .C(n6114), .D(n6113), .Y(n6974) );
  INVX12 U191 ( .A(n6979), .Y(mem_wdata[59]) );
  NOR4X2 U192 ( .A(n6120), .B(n6119), .C(n6118), .D(n6117), .Y(n6979) );
  INVX12 U193 ( .A(n7017), .Y(mem_wdata[5]) );
  NOR4X2 U194 ( .A(n6124), .B(n6123), .C(n6122), .D(n6121), .Y(n7017) );
  INVX12 U195 ( .A(n6984), .Y(mem_wdata[60]) );
  NOR4X2 U196 ( .A(n6128), .B(n6127), .C(n6126), .D(n6125), .Y(n6984) );
  INVX12 U197 ( .A(n6989), .Y(mem_wdata[61]) );
  NOR4X2 U198 ( .A(n6132), .B(n6131), .C(n6130), .D(n6129), .Y(n6989) );
  INVX12 U199 ( .A(n6999), .Y(mem_wdata[62]) );
  NOR4X2 U200 ( .A(n6136), .B(n6135), .C(n6134), .D(n6133), .Y(n6999) );
  INVX12 U201 ( .A(n7004), .Y(mem_wdata[63]) );
  NOR4X2 U202 ( .A(n6140), .B(n6139), .C(n6138), .D(n6137), .Y(n7004) );
  INVX12 U203 ( .A(n6885), .Y(mem_wdata[64]) );
  NOR4X2 U204 ( .A(n6144), .B(n6143), .C(n6142), .D(n6141), .Y(n6885) );
  INVX12 U205 ( .A(n6940), .Y(mem_wdata[65]) );
  NOR4X2 U206 ( .A(n6148), .B(n6147), .C(n6146), .D(n6145), .Y(n6940) );
  INVX12 U207 ( .A(n6995), .Y(mem_wdata[66]) );
  NOR4X2 U208 ( .A(n6152), .B(n6151), .C(n6150), .D(n6149), .Y(n6995) );
  INVX12 U209 ( .A(n7010), .Y(mem_wdata[67]) );
  NOR4X2 U210 ( .A(n6156), .B(n6155), .C(n6154), .D(n6153), .Y(n7010) );
  INVX12 U211 ( .A(n7015), .Y(mem_wdata[68]) );
  NOR4X2 U212 ( .A(n6160), .B(n6159), .C(n6158), .D(n6157), .Y(n7015) );
  INVX12 U213 ( .A(n7020), .Y(mem_wdata[69]) );
  NOR4X2 U214 ( .A(n6164), .B(n6163), .C(n6162), .D(n6161), .Y(n7020) );
  INVX12 U215 ( .A(n7022), .Y(mem_wdata[6]) );
  NOR4X2 U216 ( .A(n6168), .B(n6167), .C(n6166), .D(n6165), .Y(n7022) );
  INVX12 U217 ( .A(n7025), .Y(mem_wdata[70]) );
  NOR4X2 U218 ( .A(n6172), .B(n6171), .C(n6170), .D(n6169), .Y(n7025) );
  INVX12 U219 ( .A(n7030), .Y(mem_wdata[71]) );
  NOR4X2 U220 ( .A(n6176), .B(n6175), .C(n6174), .D(n6173), .Y(n7030) );
  INVX12 U221 ( .A(n7035), .Y(mem_wdata[72]) );
  NOR4X2 U222 ( .A(n6180), .B(n6179), .C(n6178), .D(n6177), .Y(n7035) );
  INVX12 U223 ( .A(n7044), .Y(mem_wdata[73]) );
  NOR4X2 U224 ( .A(n6184), .B(n6183), .C(n6182), .D(n6181), .Y(n7044) );
  INVX12 U225 ( .A(n6890), .Y(mem_wdata[74]) );
  NOR4X2 U226 ( .A(n6188), .B(n6187), .C(n6186), .D(n6185), .Y(n6890) );
  INVX12 U227 ( .A(n6895), .Y(mem_wdata[75]) );
  NOR4X2 U228 ( .A(n6192), .B(n6191), .C(n6190), .D(n6189), .Y(n6895) );
  INVX12 U229 ( .A(n6900), .Y(mem_wdata[76]) );
  NOR4X2 U230 ( .A(n6196), .B(n6195), .C(n6194), .D(n6193), .Y(n6900) );
  INVX12 U231 ( .A(n6905), .Y(mem_wdata[77]) );
  NOR4X2 U232 ( .A(n6200), .B(n6199), .C(n6198), .D(n6197), .Y(n6905) );
  INVX12 U233 ( .A(n6910), .Y(mem_wdata[78]) );
  NOR4X2 U234 ( .A(n6204), .B(n6203), .C(n6202), .D(n6201), .Y(n6910) );
  INVX12 U235 ( .A(n6915), .Y(mem_wdata[79]) );
  NOR4X2 U236 ( .A(n6208), .B(n6207), .C(n6206), .D(n6205), .Y(n6915) );
  INVX12 U237 ( .A(n7027), .Y(mem_wdata[7]) );
  NOR4X2 U238 ( .A(n6212), .B(n6211), .C(n6210), .D(n6209), .Y(n7027) );
  INVX12 U239 ( .A(n6920), .Y(mem_wdata[80]) );
  NOR4X2 U240 ( .A(n6216), .B(n6215), .C(n6214), .D(n6213), .Y(n6920) );
  INVX12 U241 ( .A(n6925), .Y(mem_wdata[81]) );
  NOR4X2 U242 ( .A(n6220), .B(n6219), .C(n6218), .D(n6217), .Y(n6925) );
  INVX12 U243 ( .A(n6930), .Y(mem_wdata[82]) );
  NOR4X2 U244 ( .A(n6224), .B(n6223), .C(n6222), .D(n6221), .Y(n6930) );
  INVX12 U245 ( .A(n6935), .Y(mem_wdata[83]) );
  NOR4X2 U246 ( .A(n6228), .B(n6227), .C(n6226), .D(n6225), .Y(n6935) );
  INVX12 U247 ( .A(n6945), .Y(mem_wdata[84]) );
  NOR4X2 U248 ( .A(n6232), .B(n6231), .C(n6230), .D(n6229), .Y(n6945) );
  INVX12 U249 ( .A(n6950), .Y(mem_wdata[85]) );
  NOR4X2 U250 ( .A(n6236), .B(n6235), .C(n6234), .D(n6233), .Y(n6950) );
  INVX12 U251 ( .A(n6955), .Y(mem_wdata[86]) );
  NOR4X2 U252 ( .A(n6240), .B(n6239), .C(n6238), .D(n6237), .Y(n6955) );
  INVX12 U253 ( .A(n6960), .Y(mem_wdata[87]) );
  NOR4X2 U254 ( .A(n6244), .B(n6243), .C(n6242), .D(n6241), .Y(n6960) );
  INVX12 U255 ( .A(n6965), .Y(mem_wdata[88]) );
  NOR4X2 U256 ( .A(n6248), .B(n6247), .C(n6246), .D(n6245), .Y(n6965) );
  INVX12 U257 ( .A(n6970), .Y(mem_wdata[89]) );
  NOR4X2 U258 ( .A(n6252), .B(n6251), .C(n6250), .D(n6249), .Y(n6970) );
  INVX12 U259 ( .A(n7032), .Y(mem_wdata[8]) );
  NOR4X2 U260 ( .A(n6256), .B(n6255), .C(n6254), .D(n6253), .Y(n7032) );
  INVX12 U261 ( .A(n6975), .Y(mem_wdata[90]) );
  NOR4X2 U262 ( .A(n6260), .B(n6259), .C(n6258), .D(n6257), .Y(n6975) );
  INVX12 U263 ( .A(n6980), .Y(mem_wdata[91]) );
  NOR4X2 U264 ( .A(n6264), .B(n6263), .C(n6262), .D(n6261), .Y(n6980) );
  INVX12 U265 ( .A(n6985), .Y(mem_wdata[92]) );
  NOR4X2 U266 ( .A(n6268), .B(n6267), .C(n6266), .D(n6265), .Y(n6985) );
  INVX12 U267 ( .A(n6990), .Y(mem_wdata[93]) );
  NOR4X2 U268 ( .A(n6272), .B(n6271), .C(n6270), .D(n6269), .Y(n6990) );
  INVX12 U269 ( .A(n7000), .Y(mem_wdata[94]) );
  NOR4X2 U270 ( .A(n6276), .B(n6275), .C(n6274), .D(n6273), .Y(n7000) );
  INVX12 U271 ( .A(n7005), .Y(mem_wdata[95]) );
  NOR4X2 U272 ( .A(n6280), .B(n6279), .C(n6278), .D(n6277), .Y(n7005) );
  INVX12 U273 ( .A(n6881), .Y(mem_wdata[96]) );
  NOR4X2 U274 ( .A(n6284), .B(n6283), .C(n6282), .D(n6281), .Y(n6881) );
  INVX12 U275 ( .A(n6936), .Y(mem_wdata[97]) );
  NOR4X2 U276 ( .A(n6288), .B(n6287), .C(n6286), .D(n6285), .Y(n6936) );
  INVX12 U277 ( .A(n6991), .Y(mem_wdata[98]) );
  NOR4X2 U278 ( .A(n6292), .B(n6291), .C(n6290), .D(n6289), .Y(n6991) );
  INVX12 U279 ( .A(n7006), .Y(mem_wdata[99]) );
  NOR4X2 U280 ( .A(n6296), .B(n6295), .C(n6294), .D(n6293), .Y(n7006) );
  INVX12 U281 ( .A(n7039), .Y(mem_wdata[9]) );
  NOR4X2 U282 ( .A(n6300), .B(n6299), .C(n6298), .D(n6297), .Y(n7039) );
  INVX12 U283 ( .A(n11), .Y(mem_addr[19]) );
  INVX12 U284 ( .A(n12), .Y(mem_addr[20]) );
  INVX12 U285 ( .A(n13), .Y(mem_addr[21]) );
  INVX12 U286 ( .A(n14), .Y(mem_addr[22]) );
  INVX12 U287 ( .A(n15), .Y(mem_addr[23]) );
  INVX12 U288 ( .A(n18), .Y(mem_addr[24]) );
  INVX12 U289 ( .A(n19), .Y(mem_addr[25]) );
  INVX12 U290 ( .A(n16), .Y(mem_addr[26]) );
  INVX12 U291 ( .A(n17), .Y(mem_addr[27]) );
  INVX12 U292 ( .A(n10), .Y(mem_addr[9]) );
  OA22X1 U293 ( .A0(n4003), .A1(n4411), .B0(n5708), .B1(n4004), .Y(n8290) );
  INVX12 U294 ( .A(n8290), .Y(mem_addr[18]) );
  OA22X1 U295 ( .A0(n4003), .A1(n4410), .B0(n5703), .B1(n4004), .Y(n8291) );
  INVX12 U296 ( .A(n8291), .Y(mem_addr[17]) );
  OA22X1 U297 ( .A0(n4003), .A1(n4409), .B0(n5698), .B1(n4004), .Y(n8292) );
  INVX12 U298 ( .A(n8292), .Y(mem_addr[16]) );
  OA22X1 U299 ( .A0(n4003), .A1(n4408), .B0(n5693), .B1(n9), .Y(n8293) );
  INVX12 U300 ( .A(n8293), .Y(mem_addr[15]) );
  OA22X1 U301 ( .A0(n4003), .A1(n4401), .B0(n5783), .B1(n4005), .Y(n8299) );
  INVX12 U302 ( .A(n8299), .Y(mem_addr[8]) );
  OA22X1 U303 ( .A0(n4003), .A1(n4407), .B0(n5688), .B1(n4005), .Y(n8294) );
  INVX12 U304 ( .A(n8294), .Y(mem_addr[14]) );
  OA22X1 U305 ( .A0(n4003), .A1(n4400), .B0(n5778), .B1(n9), .Y(n8300) );
  INVX12 U306 ( .A(n8300), .Y(mem_addr[7]) );
  OA22X1 U307 ( .A0(n4003), .A1(n4406), .B0(n5683), .B1(n4004), .Y(n8295) );
  INVX12 U308 ( .A(n8295), .Y(mem_addr[13]) );
  OA22X1 U309 ( .A0(n4003), .A1(n4399), .B0(n5773), .B1(n9), .Y(n8301) );
  INVX12 U310 ( .A(n8301), .Y(mem_addr[6]) );
  OA22X1 U311 ( .A0(n4003), .A1(n4405), .B0(n5678), .B1(n4005), .Y(n8296) );
  INVX12 U312 ( .A(n8296), .Y(mem_addr[12]) );
  OA22X1 U313 ( .A0(n4003), .A1(n4398), .B0(n5768), .B1(n4004), .Y(n8302) );
  INVX12 U314 ( .A(n8302), .Y(mem_addr[5]) );
  OA22X1 U315 ( .A0(n4003), .A1(n4404), .B0(n5673), .B1(n4004), .Y(n8297) );
  INVX12 U316 ( .A(n8297), .Y(mem_addr[11]) );
  OA22X1 U317 ( .A0(n4003), .A1(n4397), .B0(n5763), .B1(n4005), .Y(n8303) );
  INVX12 U318 ( .A(n8303), .Y(mem_addr[4]) );
  INVX12 U319 ( .A(n7045), .Y(mem_read) );
  OA22X1 U320 ( .A0(n4003), .A1(n4403), .B0(n5668), .B1(n4005), .Y(n8298) );
  INVX12 U321 ( .A(n8298), .Y(mem_addr[10]) );
  OA22X1 U322 ( .A0(n4003), .A1(n4396), .B0(n5758), .B1(n4005), .Y(n8304) );
  INVX12 U323 ( .A(n8304), .Y(mem_addr[3]) );
  BUFX12 U324 ( .A(n8289), .Y(mem_write) );
  CLKINVX1 U325 ( .A(n4206), .Y(n4349) );
  CLKINVX1 U326 ( .A(n6854), .Y(n4391) );
  OAI221XL U327 ( .A0(n6940), .A1(n4204), .B0(n6939), .B1(n4200), .C0(n6938), 
        .Y(proc_rdata[1]) );
  CLKINVX1 U328 ( .A(n6858), .Y(n4390) );
  CLKINVX1 U329 ( .A(n6856), .Y(n4393) );
  CLKINVX1 U330 ( .A(n6830), .Y(n4394) );
  OAI221XL U331 ( .A0(n6995), .A1(n4205), .B0(n6994), .B1(n4200), .C0(n6993), 
        .Y(proc_rdata[2]) );
  OAI221XL U332 ( .A0(n7015), .A1(n4205), .B0(n7014), .B1(n4198), .C0(n7013), 
        .Y(proc_rdata[4]) );
  OAI221XL U333 ( .A0(n7010), .A1(n4205), .B0(n7009), .B1(n4200), .C0(n7008), 
        .Y(proc_rdata[3]) );
  OAI221XL U334 ( .A0(n7030), .A1(n4205), .B0(n7029), .B1(n4198), .C0(n7028), 
        .Y(proc_rdata[7]) );
  OAI221XL U335 ( .A0(n7025), .A1(n4205), .B0(n7024), .B1(n4198), .C0(n7023), 
        .Y(proc_rdata[6]) );
  OAI221XL U336 ( .A0(n7020), .A1(n4205), .B0(n7019), .B1(n4198), .C0(n7018), 
        .Y(proc_rdata[5]) );
  OAI221XL U337 ( .A0(n7044), .A1(n4203), .B0(n7042), .B1(n4200), .C0(n7040), 
        .Y(proc_rdata[9]) );
  OAI221XL U338 ( .A0(n7035), .A1(n4205), .B0(n7034), .B1(n4199), .C0(n7033), 
        .Y(proc_rdata[8]) );
  OAI221XL U339 ( .A0(n6895), .A1(n4203), .B0(n6894), .B1(n4201), .C0(n6893), 
        .Y(proc_rdata[11]) );
  OAI221XL U340 ( .A0(n6890), .A1(n4203), .B0(n6889), .B1(n4201), .C0(n6888), 
        .Y(proc_rdata[10]) );
  OAI221XL U341 ( .A0(n6910), .A1(n4204), .B0(n6909), .B1(n4201), .C0(n6908), 
        .Y(proc_rdata[14]) );
  OAI221XL U342 ( .A0(n6905), .A1(n4204), .B0(n6904), .B1(n4201), .C0(n6903), 
        .Y(proc_rdata[13]) );
  OAI221XL U343 ( .A0(n6900), .A1(n4203), .B0(n6899), .B1(n4201), .C0(n6898), 
        .Y(proc_rdata[12]) );
  OAI221XL U344 ( .A0(n6915), .A1(n4204), .B0(n6914), .B1(n4201), .C0(n6913), 
        .Y(proc_rdata[15]) );
  OAI221XL U345 ( .A0(n7005), .A1(n4205), .B0(n7004), .B1(n4200), .C0(n7003), 
        .Y(proc_rdata[31]) );
  OAI221XL U346 ( .A0(n6990), .A1(n4205), .B0(n6989), .B1(n4200), .C0(n6988), 
        .Y(proc_rdata[29]) );
  OAI221XL U347 ( .A0(n7000), .A1(n4204), .B0(n6999), .B1(n4200), .C0(n6998), 
        .Y(proc_rdata[30]) );
  NAND3X1 U348 ( .A(n6837), .B(n4132), .C(n1333), .Y(n63) );
  NOR3X1 U349 ( .A(proc_addr[3]), .B(mem_addr[2]), .C(n4392), .Y(n6858) );
  NOR3X1 U350 ( .A(proc_addr[2]), .B(mem_addr[2]), .C(n4395), .Y(n6856) );
  NOR3X1 U351 ( .A(proc_addr[3]), .B(mem_addr[2]), .C(proc_addr[2]), .Y(n6830)
         );
  OAI22XL U352 ( .A0(n4001), .A1(n7279), .B0(n1351), .B1(n7407), .Y(n6003) );
  OAI22XL U353 ( .A0(n4000), .A1(n7311), .B0(n1350), .B1(n7439), .Y(n6143) );
  OAI22XL U354 ( .A0(n4002), .A1(n7247), .B0(n1353), .B1(n7375), .Y(n5791) );
  OAI22XL U355 ( .A0(n3997), .A1(n7248), .B0(n1352), .B1(n7376), .Y(n5947) );
  OAI22XL U356 ( .A0(n3998), .A1(n7343), .B0(n1349), .B1(n7471), .Y(n6283) );
  OAI22XL U357 ( .A0(n3998), .A1(n7344), .B0(n1349), .B1(n7472), .Y(n6287) );
  OAI22XL U358 ( .A0(n4001), .A1(n7280), .B0(n1351), .B1(n7408), .Y(n6007) );
  OAI22XL U359 ( .A0(n4001), .A1(n7281), .B0(n1351), .B1(n7409), .Y(n6011) );
  OAI22XL U360 ( .A0(n4001), .A1(n7282), .B0(n1351), .B1(n7410), .Y(n6015) );
  OAI22XL U361 ( .A0(n4000), .A1(n7312), .B0(n1350), .B1(n7440), .Y(n6147) );
  OAI22XL U362 ( .A0(n4000), .A1(n7313), .B0(n1350), .B1(n7441), .Y(n6151) );
  OAI22XL U363 ( .A0(n4000), .A1(n7314), .B0(n1350), .B1(n7442), .Y(n6155) );
  OAI22XL U364 ( .A0(n4002), .A1(n7347), .B0(n1353), .B1(n7475), .Y(n5795) );
  OAI22XL U365 ( .A0(n4001), .A1(n7249), .B0(n1351), .B1(n7377), .Y(n5991) );
  OAI22XL U366 ( .A0(n4001), .A1(n7250), .B0(n1351), .B1(n7378), .Y(n6035) );
  OAI22XL U367 ( .A0(n3997), .A1(n7251), .B0(n1351), .B1(n7379), .Y(n6079) );
  OAI22XL U368 ( .A0(n3998), .A1(n7345), .B0(n1349), .B1(n7473), .Y(n6291) );
  OAI22XL U369 ( .A0(n3998), .A1(n7346), .B0(n1349), .B1(n7474), .Y(n6295) );
  CLKINVX1 U370 ( .A(proc_addr[2]), .Y(n4392) );
  CLKINVX1 U371 ( .A(proc_addr[3]), .Y(n4395) );
  OAI22XL U372 ( .A0(n4001), .A1(n7283), .B0(n1351), .B1(n7411), .Y(n6019) );
  OAI22XL U373 ( .A0(n4001), .A1(n7284), .B0(n1351), .B1(n7412), .Y(n6023) );
  OAI22XL U374 ( .A0(n4001), .A1(n7285), .B0(n1351), .B1(n7413), .Y(n6027) );
  OAI22XL U375 ( .A0(n4001), .A1(n7286), .B0(n1351), .B1(n7414), .Y(n6031) );
  OAI22XL U376 ( .A0(n4000), .A1(n7315), .B0(n1350), .B1(n7443), .Y(n6159) );
  OAI22XL U377 ( .A0(n4000), .A1(n7316), .B0(n1350), .B1(n7444), .Y(n6163) );
  OAI22XL U378 ( .A0(n4000), .A1(n7317), .B0(n1350), .B1(n7445), .Y(n6171) );
  OAI22XL U379 ( .A0(n4000), .A1(n7318), .B0(n1350), .B1(n7446), .Y(n6175) );
  OAI22XL U380 ( .A0(n4002), .A1(n7348), .B0(n1353), .B1(n7476), .Y(n5799) );
  OAI22XL U381 ( .A0(n4002), .A1(n7349), .B0(n1353), .B1(n7477), .Y(n5803) );
  OAI22XL U382 ( .A0(n4002), .A1(n7350), .B0(n1353), .B1(n7478), .Y(n5807) );
  OAI22XL U383 ( .A0(n4000), .A1(n7252), .B0(n1350), .B1(n7380), .Y(n6123) );
  OAI22XL U384 ( .A0(n4001), .A1(n7253), .B0(n1351), .B1(n7381), .Y(n6167) );
  OAI22XL U385 ( .A0(n3999), .A1(n7254), .B0(n1348), .B1(n7382), .Y(n6211) );
  OAI22XL U386 ( .A0(n4001), .A1(n7287), .B0(n1351), .B1(n7415), .Y(n6039) );
  OAI22XL U387 ( .A0(n4001), .A1(n7288), .B0(n1351), .B1(n7416), .Y(n6043) );
  OAI22XL U388 ( .A0(n3997), .A1(n7289), .B0(n1351), .B1(n7417), .Y(n6047) );
  OAI22XL U389 ( .A0(n4000), .A1(n7319), .B0(n1350), .B1(n7447), .Y(n6179) );
  OAI22XL U390 ( .A0(n4000), .A1(n7320), .B0(n1350), .B1(n7448), .Y(n6183) );
  OAI22XL U391 ( .A0(n3999), .A1(n7321), .B0(n1350), .B1(n7449), .Y(n6187) );
  OAI22XL U392 ( .A0(n4002), .A1(n7351), .B0(n1353), .B1(n7479), .Y(n5811) );
  OAI22XL U393 ( .A0(n4002), .A1(n7352), .B0(n1353), .B1(n7480), .Y(n5815) );
  OAI22XL U394 ( .A0(n4002), .A1(n7353), .B0(n1353), .B1(n7481), .Y(n5819) );
  OAI22XL U395 ( .A0(n3999), .A1(n7255), .B0(n1348), .B1(n7383), .Y(n6255) );
  OAI22XL U396 ( .A0(n4002), .A1(n7257), .B0(n1353), .B1(n7385), .Y(n5835) );
  OAI22XL U397 ( .A0(n3998), .A1(n7256), .B0(n1349), .B1(n7384), .Y(n6299) );
  OAI22XL U398 ( .A0(n4000), .A1(n7290), .B0(n1353), .B1(n7418), .Y(n6051) );
  OAI22XL U399 ( .A0(n3995), .A1(n7291), .B0(n1347), .B1(n7419), .Y(n6055) );
  OAI22XL U400 ( .A0(n3998), .A1(n7292), .B0(n1347), .B1(n7420), .Y(n6059) );
  OAI22XL U401 ( .A0(n3999), .A1(n7322), .B0(n1352), .B1(n7450), .Y(n6191) );
  OAI22XL U402 ( .A0(n3999), .A1(n7323), .B0(n1353), .B1(n7451), .Y(n6195) );
  OAI22XL U403 ( .A0(n3999), .A1(n7324), .B0(n1349), .B1(n7452), .Y(n6199) );
  OAI22XL U404 ( .A0(n4002), .A1(n7354), .B0(n1353), .B1(n7482), .Y(n5823) );
  OAI22XL U405 ( .A0(n4002), .A1(n7355), .B0(n1353), .B1(n7483), .Y(n5827) );
  OAI22XL U406 ( .A0(n4002), .A1(n7356), .B0(n1353), .B1(n7484), .Y(n5831) );
  OAI22XL U407 ( .A0(n3997), .A1(n7258), .B0(n1348), .B1(n7386), .Y(n5879) );
  OAI22XL U408 ( .A0(n4001), .A1(n7259), .B0(n1352), .B1(n7387), .Y(n5915) );
  OAI22XL U409 ( .A0(n3996), .A1(n7260), .B0(n1352), .B1(n7388), .Y(n5919) );
  OAI22XL U410 ( .A0(n4002), .A1(n7293), .B0(n1346), .B1(n7421), .Y(n6063) );
  OAI22XL U411 ( .A0(n3997), .A1(n7294), .B0(n1346), .B1(n7422), .Y(n6067) );
  OAI22XL U412 ( .A0(n3999), .A1(n7325), .B0(n1353), .B1(n7453), .Y(n6203) );
  OAI22XL U413 ( .A0(n3999), .A1(n7326), .B0(n1348), .B1(n7454), .Y(n6207) );
  OAI22XL U414 ( .A0(n4002), .A1(n7357), .B0(n1353), .B1(n7485), .Y(n5839) );
  OAI22XL U415 ( .A0(n4002), .A1(n7358), .B0(n1353), .B1(n7486), .Y(n5843) );
  OAI22XL U416 ( .A0(n3997), .A1(n7261), .B0(n1352), .B1(n7389), .Y(n5923) );
  OAI22XL U417 ( .A0(n3995), .A1(n7262), .B0(n1352), .B1(n7390), .Y(n5927) );
  OAI22XL U418 ( .A0(n4001), .A1(n7276), .B0(n1351), .B1(n7404), .Y(n5987) );
  OAI22XL U419 ( .A0(n4001), .A1(n7277), .B0(n1351), .B1(n7405), .Y(n5995) );
  OAI22XL U420 ( .A0(n4001), .A1(n7278), .B0(n1351), .B1(n7406), .Y(n5999) );
  OAI22XL U421 ( .A0(n4000), .A1(n7308), .B0(n1350), .B1(n7436), .Y(n6131) );
  OAI22XL U422 ( .A0(n4000), .A1(n7309), .B0(n1350), .B1(n7437), .Y(n6135) );
  OAI22XL U423 ( .A0(n4000), .A1(n7310), .B0(n1350), .B1(n7438), .Y(n6139) );
  OAI22XL U424 ( .A0(n4001), .A1(n7372), .B0(n1352), .B1(n7500), .Y(n5903) );
  OAI22XL U425 ( .A0(n3996), .A1(n7373), .B0(n1346), .B1(n7501), .Y(n5907) );
  OAI22XL U426 ( .A0(n3996), .A1(n7374), .B0(n1349), .B1(n7502), .Y(n5911) );
  OAI22XL U427 ( .A0(n3998), .A1(n7340), .B0(n1349), .B1(n7468), .Y(n6271) );
  OAI22XL U428 ( .A0(n3998), .A1(n7341), .B0(n1349), .B1(n7469), .Y(n6275) );
  OAI22XL U429 ( .A0(n3998), .A1(n7342), .B0(n1349), .B1(n7470), .Y(n6279) );
  OAI22XL U430 ( .A0(n3996), .A1(n7274), .B0(n1352), .B1(n7402), .Y(n5979) );
  OAI22XL U431 ( .A0(n4001), .A1(n7275), .B0(n1351), .B1(n7403), .Y(n5983) );
  OAI22XL U432 ( .A0(n4000), .A1(n7306), .B0(n1350), .B1(n7434), .Y(n6119) );
  OAI22XL U433 ( .A0(n4000), .A1(n7307), .B0(n1350), .B1(n7435), .Y(n6127) );
  OAI22XL U434 ( .A0(n3997), .A1(n7370), .B0(n1347), .B1(n7498), .Y(n5895) );
  OAI22XL U435 ( .A0(n3996), .A1(n7371), .B0(n1351), .B1(n7499), .Y(n5899) );
  OAI22XL U436 ( .A0(n3998), .A1(n7338), .B0(n1349), .B1(n7466), .Y(n6263) );
  OAI22XL U437 ( .A0(n3998), .A1(n7339), .B0(n1349), .B1(n7467), .Y(n6267) );
  OAI22XL U438 ( .A0(n3995), .A1(n7265), .B0(n1352), .B1(n7393), .Y(n5939) );
  OAI22XL U439 ( .A0(n3998), .A1(n7266), .B0(n1352), .B1(n7394), .Y(n5943) );
  OAI22XL U440 ( .A0(n3995), .A1(n7267), .B0(n1352), .B1(n7395), .Y(n5951) );
  OAI22XL U441 ( .A0(n3997), .A1(n7268), .B0(n1352), .B1(n7396), .Y(n5955) );
  OAI22XL U442 ( .A0(n3995), .A1(n7269), .B0(n1352), .B1(n7397), .Y(n5959) );
  OAI22XL U443 ( .A0(n3996), .A1(n7270), .B0(n1352), .B1(n7398), .Y(n5963) );
  OAI22XL U444 ( .A0(n3996), .A1(n7271), .B0(n1352), .B1(n7399), .Y(n5967) );
  OAI22XL U445 ( .A0(n3996), .A1(n7272), .B0(n1352), .B1(n7400), .Y(n5971) );
  OAI22XL U446 ( .A0(n3997), .A1(n7359), .B0(n4390), .B1(n7487), .Y(n5847) );
  OAI22XL U447 ( .A0(n3997), .A1(n7360), .B0(n1348), .B1(n7488), .Y(n5851) );
  OAI22XL U448 ( .A0(n3996), .A1(n7361), .B0(n1347), .B1(n7489), .Y(n5855) );
  OAI22XL U449 ( .A0(n3997), .A1(n7362), .B0(n1348), .B1(n7490), .Y(n5859) );
  OAI22XL U450 ( .A0(n4000), .A1(n7363), .B0(n1350), .B1(n7491), .Y(n5863) );
  OAI22XL U451 ( .A0(n3995), .A1(n7364), .B0(n1352), .B1(n7492), .Y(n5867) );
  OAI22XL U452 ( .A0(n3998), .A1(n7365), .B0(n1346), .B1(n7493), .Y(n5871) );
  OAI22XL U453 ( .A0(n3995), .A1(n7366), .B0(n1347), .B1(n7494), .Y(n5875) );
  OAI22XL U454 ( .A0(n3995), .A1(n7367), .B0(n1346), .B1(n7495), .Y(n5883) );
  OAI22XL U455 ( .A0(n4002), .A1(n7368), .B0(n1347), .B1(n7496), .Y(n5887) );
  OAI22XL U456 ( .A0(n3995), .A1(n7263), .B0(n1352), .B1(n7391), .Y(n5931) );
  OAI22XL U457 ( .A0(n3997), .A1(n7264), .B0(n1352), .B1(n7392), .Y(n5935) );
  OAI22XL U458 ( .A0(n1693), .A1(n7097), .B0(n1356), .B1(n7122), .Y(n5755) );
  OAI22XL U459 ( .A0(n1695), .A1(n7098), .B0(n1359), .B1(n7123), .Y(n5760) );
  OAI22XL U460 ( .A0(n1693), .A1(n7099), .B0(n1359), .B1(n7124), .Y(n5765) );
  OAI22XL U461 ( .A0(n1693), .A1(n7100), .B0(n1354), .B1(n7125), .Y(n5770) );
  OAI22XL U462 ( .A0(n1695), .A1(n7109), .B0(n1528), .B1(n7134), .Y(n5690) );
  OAI22XL U463 ( .A0(n1693), .A1(n7110), .B0(n1356), .B1(n7135), .Y(n5695) );
  OAI22XL U464 ( .A0(n1696), .A1(n7111), .B0(n1356), .B1(n7136), .Y(n5700) );
  OAI22XL U465 ( .A0(n1696), .A1(n7112), .B0(n1358), .B1(n7137), .Y(n5705) );
  OAI22XL U466 ( .A0(n1695), .A1(n7113), .B0(n1355), .B1(n7138), .Y(n5710) );
  OAI22XL U467 ( .A0(n2628), .A1(n7114), .B0(n1354), .B1(n7139), .Y(n5715) );
  OAI22XL U468 ( .A0(n1696), .A1(n7115), .B0(n1355), .B1(n7140), .Y(n5720) );
  OAI22XL U469 ( .A0(n1701), .A1(n7116), .B0(n1356), .B1(n7141), .Y(n5725) );
  OAI22XL U470 ( .A0(n1693), .A1(n7117), .B0(n1354), .B1(n7142), .Y(n5730) );
  OAI22XL U471 ( .A0(n1696), .A1(n7118), .B0(n1356), .B1(n7143), .Y(n5735) );
  OAI22XL U472 ( .A0(n1693), .A1(n7119), .B0(n1355), .B1(n7144), .Y(n5740) );
  OAI22XL U473 ( .A0(n1696), .A1(n7120), .B0(n1580), .B1(n7145), .Y(n5745) );
  OAI22XL U474 ( .A0(n1703), .A1(n7121), .B0(n1355), .B1(n7146), .Y(n5750) );
  OAI22XL U475 ( .A0(n3999), .A1(n7047), .B0(n1348), .B1(n7072), .Y(n5754) );
  OAI22XL U476 ( .A0(n3999), .A1(n7048), .B0(n1348), .B1(n7073), .Y(n5759) );
  OAI22XL U477 ( .A0(n3999), .A1(n7049), .B0(n1352), .B1(n7074), .Y(n5764) );
  OAI22XL U478 ( .A0(n3997), .A1(n7050), .B0(n1346), .B1(n7075), .Y(n5769) );
  OAI22XL U479 ( .A0(n4002), .A1(n7051), .B0(n1353), .B1(n7076), .Y(n5774) );
  OAI22XL U480 ( .A0(n4002), .A1(n7052), .B0(n1353), .B1(n7077), .Y(n5779) );
  OAI22XL U481 ( .A0(n4002), .A1(n7053), .B0(n1353), .B1(n7078), .Y(n5784) );
  OAI22XL U482 ( .A0(n3995), .A1(n7059), .B0(n1348), .B1(n7084), .Y(n5689) );
  OAI22XL U483 ( .A0(n3997), .A1(n7060), .B0(n1347), .B1(n7085), .Y(n5694) );
  OAI22XL U484 ( .A0(n3995), .A1(n7061), .B0(n1346), .B1(n7086), .Y(n5699) );
  OAI22XL U485 ( .A0(n3996), .A1(n7062), .B0(n1346), .B1(n7087), .Y(n5704) );
  OAI22XL U486 ( .A0(n4002), .A1(n7063), .B0(n1347), .B1(n7088), .Y(n5709) );
  OAI22XL U487 ( .A0(n3997), .A1(n7064), .B0(n1351), .B1(n7089), .Y(n5714) );
  OAI22XL U488 ( .A0(n4000), .A1(n7065), .B0(n1348), .B1(n7090), .Y(n5719) );
  OAI22XL U489 ( .A0(n3995), .A1(n7066), .B0(n1347), .B1(n7091), .Y(n5724) );
  OAI22XL U490 ( .A0(n3997), .A1(n7067), .B0(n1347), .B1(n7092), .Y(n5729) );
  OAI22XL U491 ( .A0(n3995), .A1(n7068), .B0(n1346), .B1(n7093), .Y(n5734) );
  OAI22XL U492 ( .A0(n3997), .A1(n7069), .B0(n1346), .B1(n7094), .Y(n5739) );
  OAI22XL U493 ( .A0(n4001), .A1(n7070), .B0(n1347), .B1(n7095), .Y(n5744) );
  OAI22XL U494 ( .A0(n3995), .A1(n7071), .B0(n1348), .B1(n7096), .Y(n5749) );
  OAI22XL U495 ( .A0(n3998), .A1(n7054), .B0(n1349), .B1(n7079), .Y(n5664) );
  OAI22XL U496 ( .A0(n2628), .A1(n7101), .B0(n1580), .B1(n7126), .Y(n5775) );
  OAI22XL U497 ( .A0(n2628), .A1(n7102), .B0(n1580), .B1(n7127), .Y(n5780) );
  OAI22XL U498 ( .A0(n2628), .A1(n7103), .B0(n1580), .B1(n7128), .Y(n5785) );
  OAI22XL U499 ( .A0(n1697), .A1(n7104), .B0(n1356), .B1(n7129), .Y(n5665) );
  OAI22XL U500 ( .A0(n4121), .A1(n7153), .B0(n4131), .B1(n7178), .Y(n5786) );
  OAI22XL U501 ( .A0(n4393), .A1(n7105), .B0(n1357), .B1(n7130), .Y(n5670) );
  OAI22XL U502 ( .A0(n4393), .A1(n7106), .B0(n1354), .B1(n7131), .Y(n5675) );
  OAI22XL U503 ( .A0(n4393), .A1(n7107), .B0(n4391), .B1(n7132), .Y(n5680) );
  OAI22XL U504 ( .A0(n1693), .A1(n7108), .B0(n1357), .B1(n7133), .Y(n5685) );
  OAI22XL U505 ( .A0(n4394), .A1(n7055), .B0(n1347), .B1(n7080), .Y(n5669) );
  OAI22XL U506 ( .A0(n3997), .A1(n7056), .B0(n1349), .B1(n7081), .Y(n5674) );
  OAI22XL U507 ( .A0(n3996), .A1(n7057), .B0(n1348), .B1(n7082), .Y(n5679) );
  OAI22XL U508 ( .A0(n3995), .A1(n7058), .B0(n1346), .B1(n7083), .Y(n5684) );
  OAI22XL U509 ( .A0(n3996), .A1(n7273), .B0(n1352), .B1(n7401), .Y(n5975) );
  OAI22XL U510 ( .A0(n3996), .A1(n7295), .B0(n1346), .B1(n7423), .Y(n6071) );
  OAI22XL U511 ( .A0(n3995), .A1(n7296), .B0(n1347), .B1(n7424), .Y(n6075) );
  OAI22XL U512 ( .A0(n3996), .A1(n7297), .B0(n1348), .B1(n7425), .Y(n6083) );
  OAI22XL U513 ( .A0(n3995), .A1(n7298), .B0(n1347), .B1(n7426), .Y(n6087) );
  OAI22XL U514 ( .A0(n3995), .A1(n7299), .B0(n1353), .B1(n7427), .Y(n6091) );
  OAI22XL U515 ( .A0(n3995), .A1(n7300), .B0(n1348), .B1(n7428), .Y(n6095) );
  OAI22XL U516 ( .A0(n4001), .A1(n7301), .B0(n1346), .B1(n7429), .Y(n6099) );
  OAI22XL U517 ( .A0(n3997), .A1(n7302), .B0(n1346), .B1(n7430), .Y(n6103) );
  OAI22XL U518 ( .A0(n3996), .A1(n7303), .B0(n1347), .B1(n7431), .Y(n6107) );
  OAI22XL U519 ( .A0(n3997), .A1(n7304), .B0(n4390), .B1(n7432), .Y(n6111) );
  OAI22XL U520 ( .A0(n3999), .A1(n7327), .B0(n1346), .B1(n7455), .Y(n6215) );
  OAI22XL U521 ( .A0(n3999), .A1(n7328), .B0(n4390), .B1(n7456), .Y(n6219) );
  OAI22XL U522 ( .A0(n3999), .A1(n7329), .B0(n1348), .B1(n7457), .Y(n6223) );
  OAI22XL U523 ( .A0(n3999), .A1(n7330), .B0(n1348), .B1(n7458), .Y(n6227) );
  OAI22XL U524 ( .A0(n3999), .A1(n7331), .B0(n1348), .B1(n7459), .Y(n6231) );
  OAI22XL U525 ( .A0(n3999), .A1(n7332), .B0(n1348), .B1(n7460), .Y(n6235) );
  OAI22XL U526 ( .A0(n3999), .A1(n7333), .B0(n1348), .B1(n7461), .Y(n6239) );
  OAI22XL U527 ( .A0(n3999), .A1(n7334), .B0(n1348), .B1(n7462), .Y(n6243) );
  OAI22XL U528 ( .A0(n3999), .A1(n7335), .B0(n1350), .B1(n7463), .Y(n6247) );
  OAI22XL U529 ( .A0(n4394), .A1(n7369), .B0(n1347), .B1(n7497), .Y(n5891) );
  OAI22XL U530 ( .A0(n4000), .A1(n7305), .B0(n1350), .B1(n7433), .Y(n6115) );
  OAI22XL U531 ( .A0(n3998), .A1(n7336), .B0(n1349), .B1(n7464), .Y(n6251) );
  OAI22XL U532 ( .A0(n3998), .A1(n7337), .B0(n1349), .B1(n7465), .Y(n6259) );
  OAI22XL U533 ( .A0(n3998), .A1(n8281), .B0(n1349), .B1(n8282), .Y(n6835) );
  OAI21XL U534 ( .A0(proc_write), .A1(n4355), .B0(n6831), .Y(n6839) );
  CLKINVX1 U535 ( .A(proc_wdata[18]), .Y(n4374) );
  CLKINVX1 U536 ( .A(proc_wdata[19]), .Y(n4375) );
  CLKINVX1 U537 ( .A(proc_wdata[20]), .Y(n4376) );
  CLKINVX1 U538 ( .A(proc_wdata[21]), .Y(n4377) );
  CLKINVX1 U539 ( .A(proc_wdata[22]), .Y(n4378) );
  CLKINVX1 U540 ( .A(proc_wdata[23]), .Y(n4379) );
  CLKINVX1 U541 ( .A(proc_wdata[24]), .Y(n4380) );
  CLKINVX1 U542 ( .A(proc_wdata[25]), .Y(n4381) );
  CLKINVX1 U543 ( .A(proc_wdata[26]), .Y(n4382) );
  CLKINVX1 U544 ( .A(proc_wdata[27]), .Y(n4383) );
  CLKINVX1 U545 ( .A(proc_wdata[28]), .Y(n4384) );
  CLKINVX1 U546 ( .A(proc_wdata[29]), .Y(n4385) );
  CLKINVX1 U547 ( .A(proc_wdata[30]), .Y(n4386) );
  CLKINVX1 U548 ( .A(proc_wdata[31]), .Y(n4387) );
  CLKINVX1 U549 ( .A(proc_wdata[0]), .Y(n4356) );
  CLKINVX1 U550 ( .A(proc_wdata[1]), .Y(n4357) );
  CLKINVX1 U551 ( .A(proc_wdata[2]), .Y(n4358) );
  CLKINVX1 U552 ( .A(proc_wdata[3]), .Y(n4359) );
  CLKINVX1 U553 ( .A(proc_wdata[4]), .Y(n4360) );
  CLKINVX1 U554 ( .A(proc_wdata[5]), .Y(n4361) );
  CLKINVX1 U555 ( .A(proc_wdata[6]), .Y(n4362) );
  CLKINVX1 U556 ( .A(proc_wdata[7]), .Y(n4363) );
  CLKINVX1 U557 ( .A(proc_wdata[8]), .Y(n4364) );
  CLKINVX1 U558 ( .A(proc_wdata[9]), .Y(n4365) );
  CLKINVX1 U559 ( .A(proc_wdata[10]), .Y(n4366) );
  CLKINVX1 U560 ( .A(proc_wdata[11]), .Y(n4367) );
  CLKINVX1 U561 ( .A(proc_wdata[12]), .Y(n4368) );
  CLKINVX1 U562 ( .A(proc_wdata[13]), .Y(n4369) );
  CLKINVX1 U563 ( .A(proc_wdata[14]), .Y(n4370) );
  CLKINVX1 U564 ( .A(proc_wdata[15]), .Y(n4371) );
  CLKINVX1 U565 ( .A(proc_wdata[16]), .Y(n4372) );
  CLKINVX1 U566 ( .A(proc_wdata[17]), .Y(n4373) );
  CLKBUFX3 U567 ( .A(n4334), .Y(n4215) );
  CLKBUFX3 U568 ( .A(n4334), .Y(n4216) );
  CLKBUFX3 U569 ( .A(n4334), .Y(n4217) );
  CLKBUFX3 U570 ( .A(n4334), .Y(n4218) );
  CLKBUFX3 U571 ( .A(n4333), .Y(n4219) );
  CLKBUFX3 U572 ( .A(n4333), .Y(n4220) );
  CLKBUFX3 U573 ( .A(n4333), .Y(n4221) );
  CLKBUFX3 U574 ( .A(n4333), .Y(n4222) );
  CLKBUFX3 U575 ( .A(n4332), .Y(n4223) );
  CLKBUFX3 U576 ( .A(n4332), .Y(n4224) );
  CLKBUFX3 U577 ( .A(n4332), .Y(n4225) );
  CLKBUFX3 U578 ( .A(n4332), .Y(n4226) );
  CLKBUFX3 U579 ( .A(n4331), .Y(n4227) );
  CLKBUFX3 U580 ( .A(n4331), .Y(n4228) );
  CLKBUFX3 U581 ( .A(n4331), .Y(n4229) );
  CLKBUFX3 U582 ( .A(n4331), .Y(n4230) );
  CLKBUFX3 U583 ( .A(n4330), .Y(n4231) );
  CLKBUFX3 U584 ( .A(n4330), .Y(n4232) );
  CLKBUFX3 U585 ( .A(n4330), .Y(n4233) );
  CLKBUFX3 U586 ( .A(n4330), .Y(n4234) );
  CLKBUFX3 U587 ( .A(n4329), .Y(n4235) );
  CLKBUFX3 U588 ( .A(n4329), .Y(n4236) );
  CLKBUFX3 U589 ( .A(n4329), .Y(n4237) );
  CLKBUFX3 U590 ( .A(n4329), .Y(n4238) );
  CLKBUFX3 U591 ( .A(n4328), .Y(n4239) );
  CLKBUFX3 U592 ( .A(n4328), .Y(n4240) );
  CLKBUFX3 U593 ( .A(n4328), .Y(n4241) );
  CLKBUFX3 U594 ( .A(n4328), .Y(n4242) );
  CLKBUFX3 U595 ( .A(n4327), .Y(n4243) );
  CLKBUFX3 U596 ( .A(n4327), .Y(n4244) );
  CLKBUFX3 U597 ( .A(n4327), .Y(n4245) );
  CLKBUFX3 U598 ( .A(n4327), .Y(n4246) );
  CLKBUFX3 U599 ( .A(n4326), .Y(n4247) );
  CLKBUFX3 U600 ( .A(n4326), .Y(n4248) );
  CLKBUFX3 U601 ( .A(n4326), .Y(n4249) );
  CLKBUFX3 U602 ( .A(n4326), .Y(n4250) );
  CLKBUFX3 U603 ( .A(n4325), .Y(n4251) );
  CLKBUFX3 U604 ( .A(n4325), .Y(n4252) );
  CLKBUFX3 U605 ( .A(n4325), .Y(n4253) );
  CLKBUFX3 U606 ( .A(n4325), .Y(n4254) );
  CLKBUFX3 U607 ( .A(n4324), .Y(n4255) );
  CLKBUFX3 U608 ( .A(n4324), .Y(n4256) );
  CLKBUFX3 U609 ( .A(n4324), .Y(n4257) );
  CLKBUFX3 U610 ( .A(n4324), .Y(n4258) );
  CLKBUFX3 U611 ( .A(n4323), .Y(n4259) );
  CLKBUFX3 U612 ( .A(n4323), .Y(n4260) );
  CLKBUFX3 U613 ( .A(n4323), .Y(n4261) );
  CLKBUFX3 U614 ( .A(n4323), .Y(n4262) );
  CLKBUFX3 U615 ( .A(n4322), .Y(n4263) );
  CLKBUFX3 U616 ( .A(n4322), .Y(n4264) );
  CLKBUFX3 U617 ( .A(n4322), .Y(n4265) );
  CLKBUFX3 U618 ( .A(n4322), .Y(n4266) );
  CLKBUFX3 U619 ( .A(n4321), .Y(n4267) );
  CLKBUFX3 U620 ( .A(n4321), .Y(n4268) );
  CLKBUFX3 U621 ( .A(n4321), .Y(n4269) );
  CLKBUFX3 U622 ( .A(n4321), .Y(n4270) );
  CLKBUFX3 U623 ( .A(n4320), .Y(n4271) );
  CLKBUFX3 U624 ( .A(n4320), .Y(n4272) );
  CLKBUFX3 U625 ( .A(n4320), .Y(n4273) );
  CLKBUFX3 U626 ( .A(n4320), .Y(n4274) );
  CLKBUFX3 U627 ( .A(n4319), .Y(n4275) );
  CLKBUFX3 U628 ( .A(n4319), .Y(n4276) );
  CLKBUFX3 U629 ( .A(n4319), .Y(n4277) );
  CLKBUFX3 U630 ( .A(n4319), .Y(n4278) );
  CLKBUFX3 U631 ( .A(n4318), .Y(n4279) );
  CLKBUFX3 U632 ( .A(n4318), .Y(n4280) );
  CLKBUFX3 U633 ( .A(n4318), .Y(n4281) );
  CLKBUFX3 U634 ( .A(n4318), .Y(n4282) );
  CLKBUFX3 U635 ( .A(n4317), .Y(n4283) );
  CLKBUFX3 U636 ( .A(n4317), .Y(n4284) );
  CLKBUFX3 U637 ( .A(n4317), .Y(n4285) );
  CLKBUFX3 U638 ( .A(n4317), .Y(n4286) );
  CLKBUFX3 U639 ( .A(n4316), .Y(n4287) );
  CLKBUFX3 U640 ( .A(n4316), .Y(n4288) );
  CLKBUFX3 U641 ( .A(n4316), .Y(n4289) );
  CLKBUFX3 U642 ( .A(n4316), .Y(n4290) );
  CLKBUFX3 U643 ( .A(n4315), .Y(n4291) );
  CLKBUFX3 U644 ( .A(n4315), .Y(n4292) );
  CLKBUFX3 U645 ( .A(n4315), .Y(n4293) );
  CLKBUFX3 U646 ( .A(n4315), .Y(n4294) );
  CLKBUFX3 U647 ( .A(n4314), .Y(n4295) );
  CLKBUFX3 U648 ( .A(n4314), .Y(n4296) );
  CLKBUFX3 U649 ( .A(n4314), .Y(n4297) );
  CLKBUFX3 U650 ( .A(n4314), .Y(n4298) );
  CLKBUFX3 U651 ( .A(n4313), .Y(n4299) );
  CLKBUFX3 U652 ( .A(n4313), .Y(n4300) );
  CLKBUFX3 U653 ( .A(n4313), .Y(n4301) );
  CLKBUFX3 U654 ( .A(n4313), .Y(n4302) );
  CLKBUFX3 U655 ( .A(n4312), .Y(n4303) );
  CLKBUFX3 U656 ( .A(n4312), .Y(n4304) );
  CLKBUFX3 U657 ( .A(n4312), .Y(n4305) );
  CLKBUFX3 U658 ( .A(n4312), .Y(n4306) );
  CLKBUFX3 U659 ( .A(n4311), .Y(n4307) );
  CLKBUFX3 U660 ( .A(n4311), .Y(n4308) );
  CLKBUFX3 U661 ( .A(n4311), .Y(n4309) );
  CLKBUFX3 U662 ( .A(n4311), .Y(n4310) );
  CLKBUFX3 U663 ( .A(n4336), .Y(n4207) );
  CLKBUFX3 U664 ( .A(n4336), .Y(n4208) );
  CLKBUFX3 U665 ( .A(n4336), .Y(n4209) );
  CLKBUFX3 U666 ( .A(n4336), .Y(n4210) );
  CLKBUFX3 U667 ( .A(n4335), .Y(n4211) );
  CLKBUFX3 U668 ( .A(n4335), .Y(n4212) );
  CLKBUFX3 U669 ( .A(n4335), .Y(n4213) );
  CLKBUFX3 U670 ( .A(n4335), .Y(n4214) );
  CLKBUFX3 U671 ( .A(n4337), .Y(n4334) );
  CLKBUFX3 U672 ( .A(n4337), .Y(n4333) );
  CLKBUFX3 U673 ( .A(n4348), .Y(n4332) );
  CLKBUFX3 U674 ( .A(n4348), .Y(n4331) );
  CLKBUFX3 U675 ( .A(n4347), .Y(n4330) );
  CLKBUFX3 U676 ( .A(n4347), .Y(n4329) );
  CLKBUFX3 U677 ( .A(n4338), .Y(n4328) );
  CLKBUFX3 U678 ( .A(n4338), .Y(n4327) );
  CLKBUFX3 U679 ( .A(n4339), .Y(n4326) );
  CLKBUFX3 U680 ( .A(n4339), .Y(n4325) );
  CLKBUFX3 U681 ( .A(n4346), .Y(n4324) );
  CLKBUFX3 U682 ( .A(n4346), .Y(n4323) );
  CLKBUFX3 U683 ( .A(n4340), .Y(n4322) );
  CLKBUFX3 U684 ( .A(n4340), .Y(n4321) );
  CLKBUFX3 U685 ( .A(n4345), .Y(n4320) );
  CLKBUFX3 U686 ( .A(n4345), .Y(n4319) );
  CLKBUFX3 U687 ( .A(n4341), .Y(n4318) );
  CLKBUFX3 U688 ( .A(n4341), .Y(n4317) );
  CLKBUFX3 U689 ( .A(n4344), .Y(n4316) );
  CLKBUFX3 U690 ( .A(n4337), .Y(n4315) );
  CLKBUFX3 U691 ( .A(n4342), .Y(n4314) );
  CLKBUFX3 U692 ( .A(n4342), .Y(n4313) );
  CLKBUFX3 U693 ( .A(n4343), .Y(n4312) );
  CLKBUFX3 U694 ( .A(n4343), .Y(n4311) );
  CLKBUFX3 U695 ( .A(n4039), .Y(n4041) );
  CLKBUFX3 U696 ( .A(n4099), .Y(n4095) );
  CLKBUFX3 U697 ( .A(n4113), .Y(n4109) );
  CLKBUFX3 U698 ( .A(n4081), .Y(n4084) );
  CLKBUFX3 U699 ( .A(n4039), .Y(n4042) );
  CLKBUFX3 U700 ( .A(n4059), .Y(n4054) );
  CLKBUFX3 U701 ( .A(n4099), .Y(n4096) );
  CLKBUFX3 U702 ( .A(n4113), .Y(n4110) );
  CLKBUFX3 U703 ( .A(n4060), .Y(n4061) );
  CLKBUFX3 U704 ( .A(n4081), .Y(n4085) );
  CLKBUFX3 U705 ( .A(n4191), .Y(n4185) );
  CLKBUFX3 U706 ( .A(n4039), .Y(n4043) );
  CLKBUFX3 U707 ( .A(n4099), .Y(n4097) );
  CLKBUFX3 U708 ( .A(n4113), .Y(n4111) );
  CLKBUFX3 U709 ( .A(n4060), .Y(n4062) );
  CLKBUFX3 U710 ( .A(n4191), .Y(n4186) );
  CLKBUFX3 U711 ( .A(n4039), .Y(n4044) );
  CLKBUFX3 U712 ( .A(n4059), .Y(n4055) );
  CLKBUFX3 U713 ( .A(n4060), .Y(n4063) );
  CLKBUFX3 U714 ( .A(n4191), .Y(n4187) );
  CLKBUFX3 U715 ( .A(n4099), .Y(n4098) );
  CLKBUFX3 U716 ( .A(n4113), .Y(n4112) );
  CLKBUFX3 U717 ( .A(n4060), .Y(n4064) );
  CLKBUFX3 U718 ( .A(n4059), .Y(n4056) );
  CLKBUFX3 U719 ( .A(n4060), .Y(n4065) );
  CLKBUFX3 U720 ( .A(n4191), .Y(n4188) );
  CLKBUFX3 U721 ( .A(n4059), .Y(n4057) );
  CLKBUFX3 U722 ( .A(n4191), .Y(n4189) );
  CLKBUFX3 U723 ( .A(n4191), .Y(n4190) );
  CLKBUFX3 U724 ( .A(n6711), .Y(n4040) );
  CLKBUFX3 U725 ( .A(n4099), .Y(n4094) );
  CLKBUFX3 U726 ( .A(n4113), .Y(n4108) );
  CLKBUFX3 U727 ( .A(n6710), .Y(n4021) );
  CLKBUFX3 U728 ( .A(n6710), .Y(n4022) );
  CLKBUFX3 U729 ( .A(n6710), .Y(n4023) );
  CLKBUFX3 U730 ( .A(n4024), .Y(n4020) );
  CLKBUFX3 U731 ( .A(n4039), .Y(n4045) );
  CLKBUFX3 U732 ( .A(n4053), .Y(n4058) );
  INVX3 U733 ( .A(n6850), .Y(n4154) );
  INVX3 U734 ( .A(n6851), .Y(n4157) );
  INVX3 U735 ( .A(n6852), .Y(n4160) );
  INVX3 U736 ( .A(n6853), .Y(n4163) );
  INVX3 U737 ( .A(n6855), .Y(n4166) );
  CLKBUFX3 U738 ( .A(n4348), .Y(n4337) );
  CLKBUFX3 U739 ( .A(n4347), .Y(n4338) );
  CLKBUFX3 U740 ( .A(n4346), .Y(n4339) );
  CLKBUFX3 U741 ( .A(n4345), .Y(n4340) );
  CLKBUFX3 U742 ( .A(n4344), .Y(n4341) );
  CLKBUFX3 U743 ( .A(n4343), .Y(n4342) );
  CLKBUFX3 U744 ( .A(n4350), .Y(n4336) );
  CLKBUFX3 U745 ( .A(n4344), .Y(n4335) );
  CLKBUFX3 U746 ( .A(n1356), .Y(n1359) );
  CLKBUFX3 U747 ( .A(n1356), .Y(n1528) );
  CLKBUFX3 U748 ( .A(n1355), .Y(n1358) );
  CLKBUFX3 U749 ( .A(n1357), .Y(n1580) );
  INVX3 U750 ( .A(n4123), .Y(n4115) );
  INVX3 U751 ( .A(n4122), .Y(n4117) );
  INVX3 U752 ( .A(n4122), .Y(n4118) );
  INVX3 U753 ( .A(n4122), .Y(n4119) );
  INVX3 U754 ( .A(n4122), .Y(n4116) );
  INVX3 U755 ( .A(n4122), .Y(n4121) );
  INVX3 U756 ( .A(n4122), .Y(n4120) );
  CLKBUFX3 U757 ( .A(n8), .Y(n4068) );
  CLKBUFX3 U758 ( .A(n2), .Y(n4080) );
  CLKBUFX3 U759 ( .A(n2), .Y(n4079) );
  CLKBUFX3 U760 ( .A(n8), .Y(n4072) );
  CLKBUFX3 U761 ( .A(n2), .Y(n4078) );
  CLKBUFX3 U762 ( .A(n2), .Y(n4076) );
  CLKBUFX3 U763 ( .A(n8), .Y(n4070) );
  CLKBUFX3 U764 ( .A(n8), .Y(n4071) );
  CLKBUFX3 U765 ( .A(n4067), .Y(n4069) );
  CLKBUFX3 U766 ( .A(n4078), .Y(n4075) );
  CLKBUFX3 U767 ( .A(n4076), .Y(n4077) );
  CLKBUFX3 U768 ( .A(n4070), .Y(n4073) );
  CLKBUFX3 U769 ( .A(n4099), .Y(n4093) );
  CLKBUFX3 U770 ( .A(n4113), .Y(n4107) );
  CLKBUFX3 U771 ( .A(n4081), .Y(n4083) );
  CLKBUFX3 U772 ( .A(n4081), .Y(n4082) );
  CLKBUFX3 U773 ( .A(n6708), .Y(n4011) );
  CLKBUFX3 U774 ( .A(n4015), .Y(n4012) );
  CLKBUFX3 U775 ( .A(n4015), .Y(n4013) );
  CLKBUFX3 U776 ( .A(n6708), .Y(n4014) );
  CLKBUFX3 U777 ( .A(n6708), .Y(n4015) );
  CLKBUFX3 U778 ( .A(n6708), .Y(n4016) );
  CLKBUFX3 U779 ( .A(n6708), .Y(n4017) );
  CLKBUFX3 U780 ( .A(n4031), .Y(n4025) );
  CLKBUFX3 U781 ( .A(n4031), .Y(n4026) );
  CLKBUFX3 U782 ( .A(n4031), .Y(n4027) );
  CLKBUFX3 U783 ( .A(n4031), .Y(n4028) );
  CLKBUFX3 U784 ( .A(n4031), .Y(n4029) );
  CLKBUFX3 U785 ( .A(n4031), .Y(n4030) );
  CLKBUFX3 U786 ( .A(n4038), .Y(n4032) );
  CLKBUFX3 U787 ( .A(n4052), .Y(n4046) );
  CLKBUFX3 U788 ( .A(n4087), .Y(n4088) );
  CLKBUFX3 U789 ( .A(n4101), .Y(n4102) );
  CLKBUFX3 U790 ( .A(n4038), .Y(n4033) );
  CLKBUFX3 U791 ( .A(n4052), .Y(n4047) );
  CLKBUFX3 U792 ( .A(n4087), .Y(n4089) );
  CLKBUFX3 U793 ( .A(n4101), .Y(n4103) );
  CLKBUFX3 U794 ( .A(n4180), .Y(n4179) );
  CLKBUFX3 U795 ( .A(n4038), .Y(n4034) );
  CLKBUFX3 U796 ( .A(n4052), .Y(n4048) );
  CLKBUFX3 U797 ( .A(n4087), .Y(n4090) );
  CLKBUFX3 U798 ( .A(n4101), .Y(n4104) );
  CLKBUFX3 U799 ( .A(n1), .Y(n4180) );
  CLKBUFX3 U800 ( .A(n4038), .Y(n4035) );
  CLKBUFX3 U801 ( .A(n4052), .Y(n4049) );
  CLKBUFX3 U802 ( .A(n4087), .Y(n4091) );
  CLKBUFX3 U803 ( .A(n4101), .Y(n4105) );
  CLKBUFX3 U804 ( .A(n4038), .Y(n4036) );
  CLKBUFX3 U805 ( .A(n1), .Y(n4181) );
  CLKBUFX3 U806 ( .A(n4038), .Y(n4037) );
  CLKBUFX3 U807 ( .A(n4052), .Y(n4050) );
  CLKBUFX3 U808 ( .A(n4052), .Y(n4051) );
  CLKBUFX3 U809 ( .A(n1), .Y(n4182) );
  CLKBUFX3 U810 ( .A(n3), .Y(n4092) );
  CLKBUFX3 U811 ( .A(n4), .Y(n4106) );
  CLKBUFX3 U812 ( .A(n1), .Y(n4183) );
  CLKBUFX3 U813 ( .A(n1), .Y(n4184) );
  CLKBUFX3 U814 ( .A(n3), .Y(n4087) );
  CLKBUFX3 U815 ( .A(n4), .Y(n4101) );
  CLKBUFX3 U816 ( .A(n4015), .Y(n4018) );
  CLKBUFX3 U817 ( .A(n6716), .Y(n4099) );
  CLKBUFX3 U818 ( .A(n6829), .Y(n4113) );
  CLKBUFX3 U819 ( .A(n4053), .Y(n4059) );
  CLKBUFX3 U820 ( .A(n1345), .Y(n1344) );
  CLKBUFX3 U821 ( .A(n1339), .Y(n1343) );
  CLKBUFX3 U822 ( .A(n1344), .Y(n1342) );
  CLKBUFX3 U823 ( .A(n1339), .Y(n1341) );
  CLKBUFX3 U824 ( .A(n1344), .Y(n1340) );
  CLKBUFX3 U825 ( .A(mem_read), .Y(n1339) );
  CLKBUFX3 U826 ( .A(n6853), .Y(n4164) );
  INVX3 U827 ( .A(n6861), .Y(n4175) );
  INVX3 U828 ( .A(n6857), .Y(n4169) );
  INVX3 U829 ( .A(n6860), .Y(n4172) );
  CLKBUFX3 U830 ( .A(n6850), .Y(n4155) );
  CLKBUFX3 U831 ( .A(n6851), .Y(n4158) );
  CLKBUFX3 U832 ( .A(n6852), .Y(n4161) );
  CLKBUFX3 U833 ( .A(n6853), .Y(n4165) );
  CLKBUFX3 U834 ( .A(n6855), .Y(n4167) );
  CLKBUFX3 U835 ( .A(n4350), .Y(n4344) );
  CLKBUFX3 U836 ( .A(n4350), .Y(n4343) );
  CLKBUFX3 U837 ( .A(n4349), .Y(n4348) );
  CLKBUFX3 U838 ( .A(n4349), .Y(n4347) );
  CLKBUFX3 U839 ( .A(n4349), .Y(n4346) );
  CLKBUFX3 U840 ( .A(n4349), .Y(n4345) );
  CLKBUFX3 U841 ( .A(n4394), .Y(n3998) );
  CLKBUFX3 U842 ( .A(n1695), .Y(n1697) );
  CLKBUFX3 U843 ( .A(n1346), .Y(n1349) );
  CLKBUFX3 U844 ( .A(n3996), .Y(n4001) );
  CLKBUFX3 U845 ( .A(n1695), .Y(n1703) );
  CLKBUFX3 U846 ( .A(n4002), .Y(n3999) );
  CLKBUFX3 U847 ( .A(n1695), .Y(n1704) );
  CLKBUFX3 U848 ( .A(n3995), .Y(n4000) );
  CLKBUFX3 U849 ( .A(n1693), .Y(n1701) );
  CLKBUFX3 U850 ( .A(n3997), .Y(n4002) );
  CLKBUFX3 U851 ( .A(n1696), .Y(n2628) );
  CLKBUFX3 U852 ( .A(n1347), .Y(n1351) );
  CLKBUFX3 U853 ( .A(n1347), .Y(n1352) );
  CLKBUFX3 U854 ( .A(n1346), .Y(n1350) );
  CLKBUFX3 U855 ( .A(n1348), .Y(n1353) );
  INVX3 U856 ( .A(n4143), .Y(n4135) );
  INVX3 U857 ( .A(n4133), .Y(n4125) );
  INVX3 U858 ( .A(n4153), .Y(n4145) );
  INVX3 U859 ( .A(n4142), .Y(n4137) );
  INVX3 U860 ( .A(n4143), .Y(n4138) );
  INVX3 U861 ( .A(n4143), .Y(n4139) );
  INVX3 U862 ( .A(n4142), .Y(n4136) );
  INVX3 U863 ( .A(n4143), .Y(n4141) );
  INVX3 U864 ( .A(n4132), .Y(n4128) );
  INVX3 U865 ( .A(n4152), .Y(n4148) );
  INVX3 U866 ( .A(n4132), .Y(n4129) );
  INVX3 U867 ( .A(n4153), .Y(n4149) );
  INVX3 U868 ( .A(n4132), .Y(n4126) );
  INVX3 U869 ( .A(n4152), .Y(n4146) );
  INVX3 U870 ( .A(n4133), .Y(n4130) );
  INVX3 U871 ( .A(n4153), .Y(n4150) );
  INVX3 U872 ( .A(n4133), .Y(n4127) );
  INVX3 U873 ( .A(n4152), .Y(n4147) );
  INVX3 U874 ( .A(n4133), .Y(n4131) );
  INVX3 U875 ( .A(n4153), .Y(n4151) );
  CLKBUFX3 U876 ( .A(n4195), .Y(n4196) );
  CLKBUFX3 U877 ( .A(n4195), .Y(n4197) );
  CLKBUFX3 U878 ( .A(n4123), .Y(n4122) );
  CLKBUFX3 U879 ( .A(n4391), .Y(n1357) );
  CLKBUFX3 U880 ( .A(n4391), .Y(n1356) );
  CLKBUFX3 U881 ( .A(n4391), .Y(n1354) );
  CLKBUFX3 U882 ( .A(n4391), .Y(n1355) );
  INVX3 U883 ( .A(n4142), .Y(n4140) );
  INVX4 U884 ( .A(n4004), .Y(n4003) );
  CLKBUFX3 U885 ( .A(n2), .Y(n4074) );
  CLKBUFX3 U886 ( .A(n4015), .Y(n4010) );
  CLKBUFX3 U887 ( .A(n8), .Y(n4067) );
  CLKBUFX3 U888 ( .A(n4181), .Y(n4178) );
  CLKBUFX3 U889 ( .A(n3), .Y(n4086) );
  CLKBUFX3 U890 ( .A(n4), .Y(n4100) );
  CLKBUFX3 U891 ( .A(n1337), .Y(n1345) );
  CLKBUFX3 U892 ( .A(n1338), .Y(n1337) );
  CLKBUFX3 U893 ( .A(n6715), .Y(n4081) );
  CLKBUFX3 U894 ( .A(n6880), .Y(n4191) );
  CLKBUFX3 U895 ( .A(n5), .Y(n4038) );
  CLKBUFX3 U896 ( .A(n6), .Y(n4052) );
  CLKBUFX3 U897 ( .A(n7), .Y(n4031) );
  CLKBUFX3 U898 ( .A(n6860), .Y(n4173) );
  CLKBUFX3 U899 ( .A(n6687), .Y(n4008) );
  CLKBUFX3 U900 ( .A(n6620), .Y(n4006) );
  CLKBUFX3 U901 ( .A(n6654), .Y(n4007) );
  CLKBUFX3 U902 ( .A(n6706), .Y(n4009) );
  CLKBUFX3 U903 ( .A(n6861), .Y(n4176) );
  CLKBUFX3 U904 ( .A(n6857), .Y(n4170) );
  CLKBUFX3 U905 ( .A(n6860), .Y(n4174) );
  CLKBUFX3 U906 ( .A(n6850), .Y(n4156) );
  CLKBUFX3 U907 ( .A(n6851), .Y(n4159) );
  CLKBUFX3 U908 ( .A(n6852), .Y(n4162) );
  CLKBUFX3 U909 ( .A(n6855), .Y(n4168) );
  CLKINVX1 U910 ( .A(n4206), .Y(n4350) );
  CLKBUFX3 U911 ( .A(n7043), .Y(n4203) );
  CLKBUFX3 U912 ( .A(n7036), .Y(n4193) );
  CLKBUFX3 U913 ( .A(n7036), .Y(n4194) );
  CLKBUFX3 U914 ( .A(n4198), .Y(n4200) );
  CLKBUFX3 U915 ( .A(n7043), .Y(n4204) );
  CLKBUFX3 U916 ( .A(n4153), .Y(n4152) );
  CLKBUFX3 U917 ( .A(n4143), .Y(n4142) );
  CLKBUFX3 U918 ( .A(n7038), .Y(n4195) );
  CLKBUFX3 U919 ( .A(n4390), .Y(n1348) );
  CLKBUFX3 U920 ( .A(n4390), .Y(n1347) );
  CLKBUFX3 U921 ( .A(n4390), .Y(n1346) );
  CLKBUFX3 U922 ( .A(n4394), .Y(n3997) );
  CLKBUFX3 U923 ( .A(n4394), .Y(n3996) );
  CLKBUFX3 U924 ( .A(n4394), .Y(n3995) );
  CLKBUFX3 U925 ( .A(n4393), .Y(n1696) );
  CLKBUFX3 U926 ( .A(n4393), .Y(n1695) );
  CLKBUFX3 U927 ( .A(n4393), .Y(n1693) );
  CLKINVX1 U928 ( .A(n4114), .Y(n4123) );
  CLKBUFX3 U929 ( .A(n9), .Y(n4004) );
  CLKBUFX3 U930 ( .A(n9), .Y(n4005) );
  NOR2BX1 U931 ( .AN(n6717), .B(n4120), .Y(n6713) );
  NOR2BX1 U932 ( .AN(n6717), .B(n4127), .Y(n6715) );
  NOR2BX1 U933 ( .AN(n6717), .B(n4140), .Y(n6716) );
  NOR2BX1 U934 ( .AN(n6717), .B(n4151), .Y(n6829) );
  NOR2BX1 U935 ( .AN(n6717), .B(n1347), .Y(n6710) );
  CLKBUFX3 U936 ( .A(n6711), .Y(n4039) );
  NOR2BX1 U937 ( .AN(n6717), .B(n1696), .Y(n6711) );
  NOR2BX1 U938 ( .AN(n6717), .B(n4391), .Y(n6712) );
  NOR2BX1 U939 ( .AN(n6717), .B(n3999), .Y(n6880) );
  CLKINVX1 U940 ( .A(n6842), .Y(n4352) );
  CLKBUFX3 U941 ( .A(n6714), .Y(n4066) );
  CLKBUFX3 U942 ( .A(n6709), .Y(n4019) );
  INVX3 U943 ( .A(n63), .Y(n1334) );
  INVX3 U944 ( .A(n63), .Y(n1335) );
  CLKBUFX3 U945 ( .A(n4351), .Y(n1338) );
  AND3X2 U946 ( .A(n4201), .B(n4197), .C(n4205), .Y(n6687) );
  AND3X2 U947 ( .A(n4201), .B(n4194), .C(n4205), .Y(n6706) );
  AND2X2 U948 ( .A(n6622), .B(n4205), .Y(n6620) );
  AND2X2 U949 ( .A(n6622), .B(n4201), .Y(n6654) );
  AND2X2 U950 ( .A(n4193), .B(n4196), .Y(n6622) );
  CLKBUFX3 U951 ( .A(n6861), .Y(n4177) );
  CLKBUFX3 U952 ( .A(n6857), .Y(n4171) );
  AND2X2 U953 ( .A(n6859), .B(n4152), .Y(n1289) );
  CLKINVX1 U954 ( .A(n1289), .Y(n6850) );
  AND2X2 U955 ( .A(n6859), .B(n4142), .Y(n1290) );
  CLKINVX1 U956 ( .A(n1290), .Y(n6851) );
  AND2X2 U957 ( .A(n6859), .B(n4132), .Y(n1291) );
  CLKINVX1 U958 ( .A(n1291), .Y(n6852) );
  AND2X2 U959 ( .A(n6859), .B(n4123), .Y(n1292) );
  CLKINVX1 U960 ( .A(n1292), .Y(n6853) );
  AND2X2 U961 ( .A(n6859), .B(n6854), .Y(n1293) );
  CLKINVX1 U962 ( .A(n1293), .Y(n6855) );
  CLKBUFX3 U963 ( .A(n4133), .Y(n4132) );
  CLKBUFX3 U964 ( .A(proc_reset), .Y(n4206) );
  OA22X1 U965 ( .A0(n7027), .A1(n4196), .B0(n7026), .B1(n4193), .Y(n7028) );
  OA22X1 U966 ( .A0(n7022), .A1(n4196), .B0(n7021), .B1(n4193), .Y(n7023) );
  OA22X1 U967 ( .A0(n7017), .A1(n4196), .B0(n7016), .B1(n4194), .Y(n7018) );
  OA22X1 U968 ( .A0(n7012), .A1(n4196), .B0(n7011), .B1(n4193), .Y(n7013) );
  OA22X1 U969 ( .A0(n7007), .A1(n4195), .B0(n7006), .B1(n4192), .Y(n7008) );
  OA22X1 U970 ( .A0(n6992), .A1(n4197), .B0(n6991), .B1(n4194), .Y(n6993) );
  OA22X1 U971 ( .A0(n6937), .A1(n4197), .B0(n6936), .B1(n4194), .Y(n6938) );
  NOR3X1 U972 ( .A(n4392), .B(mem_addr[2]), .C(n4395), .Y(n6854) );
  NAND2X1 U973 ( .A(n4388), .B(n4389), .Y(n7038) );
  CLKBUFX3 U974 ( .A(n4202), .Y(n4205) );
  CLKBUFX3 U975 ( .A(n7043), .Y(n4202) );
  OAI221X1 U976 ( .A0(n6885), .A1(n4203), .B0(n6884), .B1(n4201), .C0(n6883), 
        .Y(proc_rdata[0]) );
  OA22X1 U977 ( .A0(n6882), .A1(n4196), .B0(n6881), .B1(n4193), .Y(n6883) );
  CLKBUFX3 U978 ( .A(n6845), .Y(n4114) );
  NAND3X1 U979 ( .A(n4392), .B(n4395), .C(mem_addr[2]), .Y(n6845) );
  CLKBUFX3 U980 ( .A(n7041), .Y(n4198) );
  CLKINVX1 U981 ( .A(n4124), .Y(n4133) );
  CLKINVX1 U982 ( .A(n4144), .Y(n4153) );
  CLKINVX1 U983 ( .A(n4134), .Y(n4143) );
  CLKBUFX3 U984 ( .A(n4199), .Y(n4201) );
  CLKBUFX3 U985 ( .A(n7041), .Y(n4199) );
  OA22X1 U986 ( .A0(n6907), .A1(n4196), .B0(n6906), .B1(n4194), .Y(n6908) );
  OA22X1 U987 ( .A0(n6902), .A1(n4196), .B0(n6901), .B1(n4193), .Y(n6903) );
  OA22X1 U988 ( .A0(n6897), .A1(n4196), .B0(n6896), .B1(n4193), .Y(n6898) );
  OA22X1 U989 ( .A0(n6892), .A1(n4196), .B0(n6891), .B1(n4193), .Y(n6893) );
  OA22X1 U990 ( .A0(n6887), .A1(n4196), .B0(n6886), .B1(n4193), .Y(n6888) );
  OA22X1 U991 ( .A0(n7039), .A1(n4196), .B0(n7037), .B1(n4193), .Y(n7040) );
  OA22X1 U992 ( .A0(n7032), .A1(n4196), .B0(n7031), .B1(n4193), .Y(n7033) );
  NOR4X1 U993 ( .A(n6432), .B(n6431), .C(n6430), .D(n6429), .Y(n6433) );
  NAND4X1 U994 ( .A(n6428), .B(n6427), .C(n6426), .D(n6425), .Y(n6429) );
  NAND4X1 U995 ( .A(n6413), .B(n6412), .C(n6411), .D(n6410), .Y(n6431) );
  NAND4X1 U996 ( .A(n6421), .B(n6420), .C(n6419), .D(n6418), .Y(n6430) );
  NOR4X1 U997 ( .A(n6399), .B(n6398), .C(n6397), .D(n6396), .Y(n6434) );
  NAND4X1 U998 ( .A(n6395), .B(n6394), .C(n6393), .D(n6392), .Y(n6396) );
  NAND4X1 U999 ( .A(n6380), .B(n6379), .C(n6378), .D(n6377), .Y(n6398) );
  NAND4X1 U1000 ( .A(n6388), .B(n6387), .C(n6386), .D(n6385), .Y(n6397) );
  NOR4X1 U1001 ( .A(n6333), .B(n6332), .C(n6331), .D(n6330), .Y(n6436) );
  NAND4X1 U1002 ( .A(n6329), .B(n6328), .C(n6327), .D(n6326), .Y(n6330) );
  NAND4X1 U1003 ( .A(n6314), .B(n6313), .C(n6312), .D(n6311), .Y(n6332) );
  NAND4X1 U1004 ( .A(n6322), .B(n6321), .C(n6320), .D(n6319), .Y(n6331) );
  NOR4X1 U1005 ( .A(n6366), .B(n6365), .C(n6364), .D(n6363), .Y(n6435) );
  NAND4X1 U1006 ( .A(n6362), .B(n6361), .C(n6360), .D(n6359), .Y(n6363) );
  NAND4X1 U1007 ( .A(n6347), .B(n6346), .C(n6345), .D(n6344), .Y(n6365) );
  NAND4X1 U1008 ( .A(n6355), .B(n6354), .C(n6353), .D(n6352), .Y(n6364) );
  AND2X2 U1009 ( .A(n6574), .B(n6573), .Y(n6838) );
  NOR4X1 U1010 ( .A(n6572), .B(n6571), .C(n6570), .D(n6569), .Y(n6573) );
  NOR4X1 U1011 ( .A(n6436), .B(n6435), .C(n6434), .D(n6433), .Y(n6574) );
  NOR4X1 U1012 ( .A(n6469), .B(n6468), .C(n6467), .D(n6466), .Y(n6572) );
  OA22X1 U1013 ( .A0(n6912), .A1(n4197), .B0(n6911), .B1(n4194), .Y(n6913) );
  CLKBUFX3 U1014 ( .A(n7036), .Y(n4192) );
  OA22X1 U1015 ( .A0(n6977), .A1(n4197), .B0(n6976), .B1(n4194), .Y(n6978) );
  OA22X1 U1016 ( .A0(n6982), .A1(n4197), .B0(n6981), .B1(n4194), .Y(n6983) );
  NOR4X1 U1017 ( .A(n6568), .B(n6567), .C(n6566), .D(n6565), .Y(n6569) );
  NAND4X1 U1018 ( .A(n6564), .B(n6563), .C(n6562), .D(n6561), .Y(n6565) );
  NAND4X1 U1019 ( .A(n6549), .B(n6548), .C(n6547), .D(n6546), .Y(n6567) );
  NAND4X1 U1020 ( .A(n6557), .B(n6556), .C(n6555), .D(n6554), .Y(n6566) );
  NOR4X1 U1021 ( .A(n6535), .B(n6534), .C(n6533), .D(n6532), .Y(n6570) );
  NAND4X1 U1022 ( .A(n6531), .B(n6530), .C(n6529), .D(n6528), .Y(n6532) );
  NAND4X1 U1023 ( .A(n6516), .B(n6515), .C(n6514), .D(n6513), .Y(n6534) );
  NAND4X1 U1024 ( .A(n6524), .B(n6523), .C(n6522), .D(n6521), .Y(n6533) );
  NOR4X1 U1025 ( .A(n6502), .B(n6501), .C(n6500), .D(n6499), .Y(n6571) );
  NAND4X1 U1026 ( .A(n6498), .B(n6497), .C(n6496), .D(n6495), .Y(n6499) );
  NAND4X1 U1027 ( .A(n6483), .B(n6482), .C(n6481), .D(n6480), .Y(n6501) );
  NAND4X1 U1028 ( .A(n6491), .B(n6490), .C(n6489), .D(n6488), .Y(n6500) );
  OA22X1 U1029 ( .A0(n7002), .A1(n4197), .B0(n7001), .B1(n4193), .Y(n7003) );
  OA22X1 U1030 ( .A0(n6997), .A1(n4197), .B0(n6996), .B1(n4194), .Y(n6998) );
  OAI21X1 U1031 ( .A0(n6832), .A1(n4421), .B0(n1336), .Y(n6842) );
  NOR2BX1 U1032 ( .AN(n6832), .B(n6838), .Y(n6708) );
  NAND2X1 U1033 ( .A(n6832), .B(n6838), .Y(n6837) );
  AND3X2 U1034 ( .A(n6837), .B(n6858), .C(n1333), .Y(n6709) );
  AND3X2 U1035 ( .A(n6837), .B(n4123), .C(n1333), .Y(n6714) );
  AND2X2 U1036 ( .A(n6837), .B(n1333), .Y(n6717) );
  CLKINVX1 U1037 ( .A(n7045), .Y(n4351) );
  OAI221XL U1038 ( .A0(n6970), .A1(n4204), .B0(n6969), .B1(n4200), .C0(n6968), 
        .Y(proc_rdata[25]) );
  OA22X1 U1039 ( .A0(n6967), .A1(n4197), .B0(n6966), .B1(n4194), .Y(n6968) );
  OAI221XL U1040 ( .A0(n6965), .A1(n4204), .B0(n6964), .B1(n4200), .C0(n6963), 
        .Y(proc_rdata[24]) );
  OA22X1 U1041 ( .A0(n6962), .A1(n4197), .B0(n6961), .B1(n4194), .Y(n6963) );
  OAI221XL U1042 ( .A0(n6960), .A1(n4204), .B0(n6959), .B1(n4200), .C0(n6958), 
        .Y(proc_rdata[23]) );
  OA22X1 U1043 ( .A0(n6957), .A1(n4197), .B0(n6956), .B1(n4194), .Y(n6958) );
  OAI221XL U1044 ( .A0(n6955), .A1(n4204), .B0(n6954), .B1(n4200), .C0(n6953), 
        .Y(proc_rdata[22]) );
  OA22X1 U1045 ( .A0(n6952), .A1(n4197), .B0(n6951), .B1(n4194), .Y(n6953) );
  OAI221XL U1046 ( .A0(n6950), .A1(n4204), .B0(n6949), .B1(n4200), .C0(n6948), 
        .Y(proc_rdata[21]) );
  OA22X1 U1047 ( .A0(n6947), .A1(n4197), .B0(n6946), .B1(n4194), .Y(n6948) );
  OAI221XL U1048 ( .A0(n6945), .A1(n4204), .B0(n6944), .B1(n4200), .C0(n6943), 
        .Y(proc_rdata[20]) );
  OA22X1 U1049 ( .A0(n6942), .A1(n4197), .B0(n6941), .B1(n4194), .Y(n6943) );
  OAI221XL U1050 ( .A0(n6935), .A1(n4204), .B0(n6934), .B1(n4200), .C0(n6933), 
        .Y(proc_rdata[19]) );
  OA22X1 U1051 ( .A0(n6932), .A1(n4197), .B0(n6931), .B1(n4194), .Y(n6933) );
  OAI221XL U1052 ( .A0(n6930), .A1(n4204), .B0(n6929), .B1(n4201), .C0(n6928), 
        .Y(proc_rdata[18]) );
  OA22X1 U1053 ( .A0(n6927), .A1(n4197), .B0(n6926), .B1(n4194), .Y(n6928) );
  OAI221XL U1054 ( .A0(n6925), .A1(n4204), .B0(n6924), .B1(n4201), .C0(n6923), 
        .Y(proc_rdata[17]) );
  OA22X1 U1055 ( .A0(n6922), .A1(n4197), .B0(n6921), .B1(n4194), .Y(n6923) );
  OAI221XL U1056 ( .A0(n6920), .A1(n4203), .B0(n6919), .B1(n4201), .C0(n6918), 
        .Y(proc_rdata[16]) );
  OA22X1 U1057 ( .A0(n6917), .A1(n4197), .B0(n6916), .B1(n4193), .Y(n6918) );
  OA22X1 U1058 ( .A0(n6987), .A1(n4197), .B0(n6986), .B1(n4194), .Y(n6988) );
  INVX3 U1059 ( .A(n1309), .Y(n4397) );
  INVX3 U1060 ( .A(n1310), .Y(n4398) );
  INVX3 U1061 ( .A(n1311), .Y(n4399) );
  INVX3 U1062 ( .A(n1312), .Y(n4400) );
  INVX3 U1063 ( .A(n1313), .Y(n4401) );
  INVX3 U1064 ( .A(n1314), .Y(n4402) );
  INVX3 U1065 ( .A(n1315), .Y(n4403) );
  INVX3 U1066 ( .A(n1316), .Y(n4404) );
  INVX3 U1067 ( .A(n1317), .Y(n4405) );
  INVX3 U1068 ( .A(n1318), .Y(n4406) );
  INVX3 U1069 ( .A(n1319), .Y(n4407) );
  INVX3 U1070 ( .A(n1320), .Y(n4408) );
  INVX3 U1071 ( .A(n1321), .Y(n4409) );
  INVX3 U1072 ( .A(n1322), .Y(n4410) );
  INVX3 U1073 ( .A(n1323), .Y(n4411) );
  INVX3 U1074 ( .A(n1324), .Y(n4412) );
  INVX3 U1075 ( .A(n1325), .Y(n4413) );
  INVX3 U1076 ( .A(n1326), .Y(n4414) );
  INVX3 U1077 ( .A(n1327), .Y(n4415) );
  INVX3 U1078 ( .A(n1328), .Y(n4416) );
  INVX3 U1079 ( .A(n1329), .Y(n4417) );
  INVX3 U1080 ( .A(n1330), .Y(n4418) );
  INVX3 U1081 ( .A(n1331), .Y(n4419) );
  INVX3 U1082 ( .A(n1308), .Y(n4396) );
  INVX3 U1083 ( .A(n1332), .Y(n4420) );
  NOR2X2 U1084 ( .A(n4421), .B(n7045), .Y(n6859) );
  AND2X2 U1085 ( .A(n6859), .B(n6858), .Y(n1294) );
  CLKINVX1 U1086 ( .A(n1294), .Y(n6860) );
  AND2X2 U1087 ( .A(n6859), .B(n6830), .Y(n1295) );
  CLKINVX1 U1088 ( .A(n1295), .Y(n6861) );
  AND2X2 U1089 ( .A(n6859), .B(n6856), .Y(n1296) );
  CLKINVX1 U1090 ( .A(n1296), .Y(n6857) );
  BUFX16 U1091 ( .A(proc_addr[4]), .Y(mem_addr[2]) );
  OAI22XL U1092 ( .A0(n1703), .A1(n7535), .B0(n1359), .B1(n7663), .Y(n6004) );
  OAI22XL U1093 ( .A0(n4138), .A1(n8047), .B0(n4149), .B1(n8175), .Y(n6002) );
  OAI22XL U1094 ( .A0(n4118), .A1(n7791), .B0(n4129), .B1(n7919), .Y(n6001) );
  OAI22XL U1095 ( .A0(n1703), .A1(n7536), .B0(n1359), .B1(n7664), .Y(n6008) );
  OAI22XL U1096 ( .A0(n4138), .A1(n8048), .B0(n4149), .B1(n8176), .Y(n6006) );
  OAI22XL U1097 ( .A0(n4118), .A1(n7792), .B0(n4129), .B1(n7920), .Y(n6005) );
  OAI22XL U1098 ( .A0(n1703), .A1(n7537), .B0(n1359), .B1(n7665), .Y(n6012) );
  OAI22XL U1099 ( .A0(n4138), .A1(n8049), .B0(n4149), .B1(n8177), .Y(n6010) );
  OAI22XL U1100 ( .A0(n4118), .A1(n7793), .B0(n4129), .B1(n7921), .Y(n6009) );
  OAI22XL U1101 ( .A0(n1703), .A1(n7538), .B0(n1359), .B1(n7666), .Y(n6016) );
  OAI22XL U1102 ( .A0(n4138), .A1(n8050), .B0(n4149), .B1(n8178), .Y(n6014) );
  OAI22XL U1103 ( .A0(n4118), .A1(n7794), .B0(n4129), .B1(n7922), .Y(n6013) );
  OAI22XL U1104 ( .A0(n1703), .A1(n7539), .B0(n1359), .B1(n7667), .Y(n6020) );
  OAI22XL U1105 ( .A0(n4138), .A1(n8051), .B0(n4149), .B1(n8179), .Y(n6018) );
  OAI22XL U1106 ( .A0(n4118), .A1(n7795), .B0(n4129), .B1(n7923), .Y(n6017) );
  OAI22XL U1107 ( .A0(n1703), .A1(n7540), .B0(n1359), .B1(n7668), .Y(n6024) );
  OAI22XL U1108 ( .A0(n4138), .A1(n8052), .B0(n4149), .B1(n8180), .Y(n6022) );
  OAI22XL U1109 ( .A0(n4118), .A1(n7796), .B0(n4129), .B1(n7924), .Y(n6021) );
  OAI22XL U1110 ( .A0(n1703), .A1(n7541), .B0(n1359), .B1(n7669), .Y(n6028) );
  OAI22XL U1111 ( .A0(n4138), .A1(n8053), .B0(n4149), .B1(n8181), .Y(n6026) );
  OAI22XL U1112 ( .A0(n4118), .A1(n7797), .B0(n4129), .B1(n7925), .Y(n6025) );
  OAI22XL U1113 ( .A0(n1701), .A1(n7567), .B0(n1358), .B1(n7695), .Y(n6144) );
  OAI22XL U1114 ( .A0(n4136), .A1(n8079), .B0(n4147), .B1(n8207), .Y(n6142) );
  OAI22XL U1115 ( .A0(n4116), .A1(n7823), .B0(n4127), .B1(n7951), .Y(n6141) );
  OAI22XL U1116 ( .A0(n1701), .A1(n7568), .B0(n1358), .B1(n7696), .Y(n6148) );
  OAI22XL U1117 ( .A0(n4136), .A1(n8080), .B0(n4147), .B1(n8208), .Y(n6146) );
  OAI22XL U1118 ( .A0(n4116), .A1(n7824), .B0(n4127), .B1(n7952), .Y(n6145) );
  OAI22XL U1119 ( .A0(n1701), .A1(n7569), .B0(n1358), .B1(n7697), .Y(n6152) );
  OAI22XL U1120 ( .A0(n4136), .A1(n8081), .B0(n4147), .B1(n8209), .Y(n6150) );
  OAI22XL U1121 ( .A0(n4116), .A1(n7825), .B0(n4127), .B1(n7953), .Y(n6149) );
  OAI22XL U1122 ( .A0(n1701), .A1(n7570), .B0(n1358), .B1(n7698), .Y(n6156) );
  OAI22XL U1123 ( .A0(n4136), .A1(n8082), .B0(n4147), .B1(n8210), .Y(n6154) );
  OAI22XL U1124 ( .A0(n4116), .A1(n7826), .B0(n4127), .B1(n7954), .Y(n6153) );
  OAI22XL U1125 ( .A0(n1701), .A1(n7571), .B0(n1358), .B1(n7699), .Y(n6160) );
  OAI22XL U1126 ( .A0(n4136), .A1(n8083), .B0(n4147), .B1(n8211), .Y(n6158) );
  OAI22XL U1127 ( .A0(n4116), .A1(n7827), .B0(n4127), .B1(n7955), .Y(n6157) );
  OAI22XL U1128 ( .A0(n1701), .A1(n7572), .B0(n1358), .B1(n7700), .Y(n6164) );
  OAI22XL U1129 ( .A0(n4136), .A1(n8084), .B0(n4147), .B1(n8212), .Y(n6162) );
  OAI22XL U1130 ( .A0(n4116), .A1(n7828), .B0(n4127), .B1(n7956), .Y(n6161) );
  OAI22XL U1131 ( .A0(n1701), .A1(n7573), .B0(n1358), .B1(n7701), .Y(n6172) );
  OAI22XL U1132 ( .A0(n4136), .A1(n8085), .B0(n4147), .B1(n8213), .Y(n6170) );
  OAI22XL U1133 ( .A0(n4116), .A1(n7829), .B0(n4127), .B1(n7957), .Y(n6169) );
  OAI22XL U1134 ( .A0(n1697), .A1(n7599), .B0(n1354), .B1(n7727), .Y(n6284) );
  OAI22XL U1135 ( .A0(n4135), .A1(n8111), .B0(n4145), .B1(n8239), .Y(n6282) );
  OAI22XL U1136 ( .A0(n4115), .A1(n7855), .B0(n4125), .B1(n7983), .Y(n6281) );
  OAI22XL U1137 ( .A0(n1697), .A1(n7600), .B0(n1354), .B1(n7728), .Y(n6288) );
  OAI22XL U1138 ( .A0(n4135), .A1(n8112), .B0(n4145), .B1(n8240), .Y(n6286) );
  OAI22XL U1139 ( .A0(n4115), .A1(n7856), .B0(n4125), .B1(n7984), .Y(n6285) );
  OAI22XL U1140 ( .A0(n1697), .A1(n7601), .B0(n1354), .B1(n7729), .Y(n6292) );
  OAI22XL U1141 ( .A0(n4135), .A1(n8113), .B0(n4145), .B1(n8241), .Y(n6290) );
  OAI22XL U1142 ( .A0(n4115), .A1(n7857), .B0(n4125), .B1(n7985), .Y(n6289) );
  OAI22XL U1143 ( .A0(n1697), .A1(n7602), .B0(n1354), .B1(n7730), .Y(n6296) );
  OAI22XL U1144 ( .A0(n4135), .A1(n8114), .B0(n4145), .B1(n8242), .Y(n6294) );
  OAI22XL U1145 ( .A0(n4115), .A1(n7858), .B0(n4125), .B1(n7986), .Y(n6293) );
  OAI22XL U1146 ( .A0(n2628), .A1(n7603), .B0(n1580), .B1(n7731), .Y(n5796) );
  OAI22XL U1147 ( .A0(n4141), .A1(n8115), .B0(n4151), .B1(n8243), .Y(n5794) );
  OAI22XL U1148 ( .A0(n4121), .A1(n7859), .B0(n4131), .B1(n7987), .Y(n5793) );
  OAI22XL U1149 ( .A0(n2628), .A1(n7604), .B0(n1580), .B1(n7732), .Y(n5800) );
  OAI22XL U1150 ( .A0(n4141), .A1(n8116), .B0(n4151), .B1(n8244), .Y(n5798) );
  OAI22XL U1151 ( .A0(n4121), .A1(n7860), .B0(n4131), .B1(n7988), .Y(n5797) );
  OAI22XL U1152 ( .A0(n2628), .A1(n7605), .B0(n1580), .B1(n7733), .Y(n5804) );
  OAI22XL U1153 ( .A0(n4141), .A1(n8117), .B0(n4151), .B1(n8245), .Y(n5802) );
  OAI22XL U1154 ( .A0(n4121), .A1(n7861), .B0(n4131), .B1(n7989), .Y(n5801) );
  OAI22XL U1155 ( .A0(n2628), .A1(n7606), .B0(n1580), .B1(n7734), .Y(n5808) );
  OAI22XL U1156 ( .A0(n4141), .A1(n8118), .B0(n4151), .B1(n8246), .Y(n5806) );
  OAI22XL U1157 ( .A0(n4121), .A1(n7862), .B0(n4131), .B1(n7990), .Y(n5805) );
  OAI22XL U1158 ( .A0(n2628), .A1(n7503), .B0(n1580), .B1(n7631), .Y(n5792) );
  OAI22XL U1159 ( .A0(n4141), .A1(n8015), .B0(n4151), .B1(n8143), .Y(n5790) );
  OAI22XL U1160 ( .A0(n4121), .A1(n7759), .B0(n4131), .B1(n7887), .Y(n5789) );
  OAI22XL U1161 ( .A0(n1704), .A1(n7504), .B0(n1528), .B1(n7632), .Y(n5948) );
  OAI22XL U1162 ( .A0(n4139), .A1(n8016), .B0(n4150), .B1(n8144), .Y(n5946) );
  OAI22XL U1163 ( .A0(n4119), .A1(n7760), .B0(n4130), .B1(n7888), .Y(n5945) );
  OAI22XL U1164 ( .A0(n1703), .A1(n7505), .B0(n1359), .B1(n7633), .Y(n5992) );
  OAI22XL U1165 ( .A0(n4138), .A1(n8017), .B0(n4149), .B1(n8145), .Y(n5990) );
  OAI22XL U1166 ( .A0(n4118), .A1(n7761), .B0(n4129), .B1(n7889), .Y(n5989) );
  OAI22XL U1167 ( .A0(n1703), .A1(n7506), .B0(n1359), .B1(n7634), .Y(n6036) );
  OAI22XL U1168 ( .A0(n4138), .A1(n8018), .B0(n4149), .B1(n8146), .Y(n6034) );
  OAI22XL U1169 ( .A0(n4118), .A1(n7762), .B0(n4129), .B1(n7890), .Y(n6033) );
  OAI22XL U1170 ( .A0(n1696), .A1(n7507), .B0(n1358), .B1(n7635), .Y(n6080) );
  OAI22XL U1171 ( .A0(n4137), .A1(n8019), .B0(n4148), .B1(n8147), .Y(n6078) );
  OAI22XL U1172 ( .A0(n4117), .A1(n7763), .B0(n4128), .B1(n7891), .Y(n6077) );
  OAI22XL U1173 ( .A0(n1701), .A1(n7508), .B0(n1358), .B1(n7636), .Y(n6124) );
  OAI22XL U1174 ( .A0(n4136), .A1(n8020), .B0(n4147), .B1(n8148), .Y(n6122) );
  OAI22XL U1175 ( .A0(n4116), .A1(n7764), .B0(n4127), .B1(n7892), .Y(n6121) );
  OAI22XL U1176 ( .A0(n1703), .A1(n7509), .B0(n1359), .B1(n7637), .Y(n6168) );
  OAI22XL U1177 ( .A0(n4138), .A1(n8021), .B0(n4149), .B1(n8149), .Y(n6166) );
  OAI22XL U1178 ( .A0(n4118), .A1(n7765), .B0(n4129), .B1(n7893), .Y(n6165) );
  OAI22XL U1179 ( .A0(n1704), .A1(n7510), .B0(n1357), .B1(n7638), .Y(n6212) );
  OAI22XL U1180 ( .A0(n4140), .A1(n8022), .B0(n4146), .B1(n8150), .Y(n6210) );
  OAI22XL U1181 ( .A0(n4120), .A1(n7766), .B0(n4126), .B1(n7894), .Y(n6209) );
  NAND2X1 U1182 ( .A(proc_addr_1), .B(proc_addr_0), .Y(n7036) );
  NAND2X1 U1183 ( .A(proc_addr_1), .B(n4388), .Y(n7043) );
  NAND2X1 U1184 ( .A(proc_addr_0), .B(n4389), .Y(n7041) );
  OAI221XL U1185 ( .A0(n6975), .A1(n4204), .B0(n6974), .B1(n4200), .C0(n6973), 
        .Y(proc_rdata[26]) );
  OA22X1 U1186 ( .A0(n6972), .A1(n4197), .B0(n6971), .B1(n4194), .Y(n6973) );
  CLKINVX1 U1187 ( .A(proc_addr_0), .Y(n4388) );
  CLKINVX1 U1188 ( .A(proc_addr_1), .Y(n4389) );
  NAND3X1 U1189 ( .A(n7046), .B(n8272), .C(n7045), .Y(proc_stall) );
  CLKBUFX3 U1190 ( .A(n6846), .Y(n4124) );
  NAND3X1 U1191 ( .A(proc_addr[2]), .B(n4395), .C(mem_addr[2]), .Y(n6846) );
  CLKBUFX3 U1192 ( .A(n6849), .Y(n4144) );
  NAND3X1 U1193 ( .A(proc_addr[3]), .B(proc_addr[2]), .C(mem_addr[2]), .Y(
        n6849) );
  CLKBUFX3 U1194 ( .A(n6847), .Y(n4134) );
  NAND3X1 U1195 ( .A(proc_addr[3]), .B(n4392), .C(mem_addr[2]), .Y(n6847) );
  OAI22XL U1196 ( .A0(n1703), .A1(n7542), .B0(n1359), .B1(n7670), .Y(n6032) );
  OAI22XL U1197 ( .A0(n4138), .A1(n8054), .B0(n4149), .B1(n8182), .Y(n6030) );
  OAI22XL U1198 ( .A0(n4118), .A1(n7798), .B0(n4129), .B1(n7926), .Y(n6029) );
  OAI22XL U1199 ( .A0(n1703), .A1(n7543), .B0(n1359), .B1(n7671), .Y(n6040) );
  OAI22XL U1200 ( .A0(n4138), .A1(n8055), .B0(n4149), .B1(n8183), .Y(n6038) );
  OAI22XL U1201 ( .A0(n4118), .A1(n7799), .B0(n4129), .B1(n7927), .Y(n6037) );
  OAI22XL U1202 ( .A0(n1703), .A1(n7544), .B0(n1359), .B1(n7672), .Y(n6044) );
  OAI22XL U1203 ( .A0(n4138), .A1(n8056), .B0(n4149), .B1(n8184), .Y(n6042) );
  OAI22XL U1204 ( .A0(n4118), .A1(n7800), .B0(n4129), .B1(n7928), .Y(n6041) );
  OAI22XL U1205 ( .A0(n1696), .A1(n7545), .B0(n1355), .B1(n7673), .Y(n6048) );
  OAI22XL U1206 ( .A0(n4137), .A1(n8057), .B0(n4148), .B1(n8185), .Y(n6046) );
  OAI22XL U1207 ( .A0(n4117), .A1(n7801), .B0(n4128), .B1(n7929), .Y(n6045) );
  OAI22XL U1208 ( .A0(n1696), .A1(n7546), .B0(n1357), .B1(n7674), .Y(n6052) );
  OAI22XL U1209 ( .A0(n4137), .A1(n8058), .B0(n4148), .B1(n8186), .Y(n6050) );
  OAI22XL U1210 ( .A0(n4117), .A1(n7802), .B0(n4128), .B1(n7930), .Y(n6049) );
  OAI22XL U1211 ( .A0(n1696), .A1(n7547), .B0(n1354), .B1(n7675), .Y(n6056) );
  OAI22XL U1212 ( .A0(n4137), .A1(n8059), .B0(n4148), .B1(n8187), .Y(n6054) );
  OAI22XL U1213 ( .A0(n4117), .A1(n7803), .B0(n4128), .B1(n7931), .Y(n6053) );
  OAI22XL U1214 ( .A0(n4137), .A1(n8060), .B0(n4148), .B1(n8188), .Y(n6058) );
  OAI22XL U1215 ( .A0(n1701), .A1(n7548), .B0(n1359), .B1(n7676), .Y(n6060) );
  OAI22XL U1216 ( .A0(n4117), .A1(n7804), .B0(n4128), .B1(n7932), .Y(n6057) );
  OAI22XL U1217 ( .A0(n4137), .A1(n8061), .B0(n4148), .B1(n8189), .Y(n6062) );
  OAI22XL U1218 ( .A0(n4117), .A1(n7805), .B0(n4128), .B1(n7933), .Y(n6061) );
  OAI22XL U1219 ( .A0(n1693), .A1(n7549), .B0(n1355), .B1(n7677), .Y(n6064) );
  OAI22XL U1220 ( .A0(n4137), .A1(n8062), .B0(n4148), .B1(n8190), .Y(n6066) );
  OAI22XL U1221 ( .A0(n4117), .A1(n7806), .B0(n4128), .B1(n7934), .Y(n6065) );
  OAI22XL U1222 ( .A0(n1704), .A1(n7550), .B0(n1357), .B1(n7678), .Y(n6068) );
  OAI22XL U1223 ( .A0(n1701), .A1(n7574), .B0(n1358), .B1(n7702), .Y(n6176) );
  OAI22XL U1224 ( .A0(n4136), .A1(n8086), .B0(n4147), .B1(n8214), .Y(n6174) );
  OAI22XL U1225 ( .A0(n4116), .A1(n7830), .B0(n4127), .B1(n7958), .Y(n6173) );
  OAI22XL U1226 ( .A0(n1701), .A1(n7575), .B0(n1358), .B1(n7703), .Y(n6180) );
  OAI22XL U1227 ( .A0(n4136), .A1(n8087), .B0(n4147), .B1(n8215), .Y(n6178) );
  OAI22XL U1228 ( .A0(n4116), .A1(n7831), .B0(n4127), .B1(n7959), .Y(n6177) );
  OAI22XL U1229 ( .A0(n1701), .A1(n7576), .B0(n1358), .B1(n7704), .Y(n6184) );
  OAI22XL U1230 ( .A0(n4136), .A1(n8088), .B0(n4147), .B1(n8216), .Y(n6182) );
  OAI22XL U1231 ( .A0(n4116), .A1(n7832), .B0(n4127), .B1(n7960), .Y(n6181) );
  OAI22XL U1232 ( .A0(n1696), .A1(n7577), .B0(n1355), .B1(n7705), .Y(n6188) );
  OAI22XL U1233 ( .A0(n4140), .A1(n8089), .B0(n4146), .B1(n8217), .Y(n6186) );
  OAI22XL U1234 ( .A0(n4120), .A1(n7833), .B0(n4126), .B1(n7961), .Y(n6185) );
  OAI22XL U1235 ( .A0(n1697), .A1(n7578), .B0(n1528), .B1(n7706), .Y(n6192) );
  OAI22XL U1236 ( .A0(n4137), .A1(n8090), .B0(n4146), .B1(n8218), .Y(n6190) );
  OAI22XL U1237 ( .A0(n4117), .A1(n7834), .B0(n4126), .B1(n7962), .Y(n6189) );
  OAI22XL U1238 ( .A0(n1695), .A1(n7579), .B0(n1354), .B1(n7707), .Y(n6196) );
  OAI22XL U1239 ( .A0(n4137), .A1(n8091), .B0(n4146), .B1(n8219), .Y(n6194) );
  OAI22XL U1240 ( .A0(n4117), .A1(n7835), .B0(n4126), .B1(n7963), .Y(n6193) );
  OAI22XL U1241 ( .A0(n1693), .A1(n7580), .B0(n1356), .B1(n7708), .Y(n6200) );
  OAI22XL U1242 ( .A0(n4137), .A1(n8092), .B0(n4146), .B1(n8220), .Y(n6198) );
  OAI22XL U1243 ( .A0(n4117), .A1(n7836), .B0(n4126), .B1(n7964), .Y(n6197) );
  OAI22XL U1244 ( .A0(n1696), .A1(n7581), .B0(n1580), .B1(n7709), .Y(n6204) );
  OAI22XL U1245 ( .A0(n4137), .A1(n8093), .B0(n4146), .B1(n8221), .Y(n6202) );
  OAI22XL U1246 ( .A0(n4117), .A1(n7837), .B0(n4126), .B1(n7965), .Y(n6201) );
  OAI22XL U1247 ( .A0(n2628), .A1(n7607), .B0(n1580), .B1(n7735), .Y(n5812) );
  OAI22XL U1248 ( .A0(n4141), .A1(n8119), .B0(n4151), .B1(n8247), .Y(n5810) );
  OAI22XL U1249 ( .A0(n4121), .A1(n7863), .B0(n4131), .B1(n7991), .Y(n5809) );
  OAI22XL U1250 ( .A0(n2628), .A1(n7608), .B0(n1580), .B1(n7736), .Y(n5816) );
  OAI22XL U1251 ( .A0(n4141), .A1(n8120), .B0(n4151), .B1(n8248), .Y(n5814) );
  OAI22XL U1252 ( .A0(n4121), .A1(n7864), .B0(n4131), .B1(n7992), .Y(n5813) );
  OAI22XL U1253 ( .A0(n2628), .A1(n7609), .B0(n1580), .B1(n7737), .Y(n5820) );
  OAI22XL U1254 ( .A0(n4141), .A1(n8121), .B0(n4151), .B1(n8249), .Y(n5818) );
  OAI22XL U1255 ( .A0(n4121), .A1(n7865), .B0(n4131), .B1(n7993), .Y(n5817) );
  OAI22XL U1256 ( .A0(n2628), .A1(n7610), .B0(n1580), .B1(n7738), .Y(n5824) );
  OAI22XL U1257 ( .A0(n4141), .A1(n8122), .B0(n4151), .B1(n8250), .Y(n5822) );
  OAI22XL U1258 ( .A0(n4121), .A1(n7866), .B0(n4131), .B1(n7994), .Y(n5821) );
  OAI22XL U1259 ( .A0(n2628), .A1(n7611), .B0(n1580), .B1(n7739), .Y(n5828) );
  OAI22XL U1260 ( .A0(n4141), .A1(n8123), .B0(n4151), .B1(n8251), .Y(n5826) );
  OAI22XL U1261 ( .A0(n4121), .A1(n7867), .B0(n4131), .B1(n7995), .Y(n5825) );
  OAI22XL U1262 ( .A0(n2628), .A1(n7612), .B0(n1580), .B1(n7740), .Y(n5832) );
  OAI22XL U1263 ( .A0(n4141), .A1(n8124), .B0(n4151), .B1(n8252), .Y(n5830) );
  OAI22XL U1264 ( .A0(n4121), .A1(n7868), .B0(n4131), .B1(n7996), .Y(n5829) );
  OAI22XL U1265 ( .A0(n2628), .A1(n7613), .B0(n1580), .B1(n7741), .Y(n5840) );
  OAI22XL U1266 ( .A0(n4141), .A1(n8125), .B0(n4151), .B1(n8253), .Y(n5838) );
  OAI22XL U1267 ( .A0(n4121), .A1(n7869), .B0(n4131), .B1(n7997), .Y(n5837) );
  OAI22XL U1268 ( .A0(n2628), .A1(n7614), .B0(n1580), .B1(n7742), .Y(n5844) );
  OAI22XL U1269 ( .A0(n4141), .A1(n8126), .B0(n4151), .B1(n8254), .Y(n5842) );
  OAI22XL U1270 ( .A0(n4121), .A1(n7870), .B0(n4131), .B1(n7998), .Y(n5841) );
  OAI22XL U1271 ( .A0(n2628), .A1(n7511), .B0(n1357), .B1(n7639), .Y(n6256) );
  OAI22XL U1272 ( .A0(n4140), .A1(n8023), .B0(n4146), .B1(n8151), .Y(n6254) );
  OAI22XL U1273 ( .A0(n4120), .A1(n7767), .B0(n4126), .B1(n7895), .Y(n6253) );
  OAI22XL U1274 ( .A0(n1697), .A1(n7512), .B0(n1354), .B1(n7640), .Y(n6300) );
  OAI22XL U1275 ( .A0(n4135), .A1(n8024), .B0(n4145), .B1(n8152), .Y(n6298) );
  OAI22XL U1276 ( .A0(n4115), .A1(n7768), .B0(n4125), .B1(n7896), .Y(n6297) );
  OAI22XL U1277 ( .A0(n2628), .A1(n7513), .B0(n1580), .B1(n7641), .Y(n5836) );
  OAI22XL U1278 ( .A0(n4141), .A1(n8025), .B0(n4151), .B1(n8153), .Y(n5834) );
  OAI22XL U1279 ( .A0(n4121), .A1(n7769), .B0(n4131), .B1(n7897), .Y(n5833) );
  OAI22XL U1280 ( .A0(n1703), .A1(n7514), .B0(n1357), .B1(n7642), .Y(n5880) );
  OAI22XL U1281 ( .A0(n4140), .A1(n8026), .B0(n4147), .B1(n8154), .Y(n5878) );
  OAI22XL U1282 ( .A0(n4120), .A1(n7770), .B0(n4131), .B1(n7898), .Y(n5877) );
  OAI22XL U1283 ( .A0(n1704), .A1(n7515), .B0(n1528), .B1(n7643), .Y(n5916) );
  OAI22XL U1284 ( .A0(n4139), .A1(n8027), .B0(n4150), .B1(n8155), .Y(n5914) );
  OAI22XL U1285 ( .A0(n4119), .A1(n7771), .B0(n4130), .B1(n7899), .Y(n5913) );
  OAI22XL U1286 ( .A0(n1704), .A1(n7516), .B0(n1528), .B1(n7644), .Y(n5920) );
  OAI22XL U1287 ( .A0(n4139), .A1(n8028), .B0(n4150), .B1(n8156), .Y(n5918) );
  OAI22XL U1288 ( .A0(n4119), .A1(n7772), .B0(n4130), .B1(n7900), .Y(n5917) );
  OAI22XL U1289 ( .A0(n1704), .A1(n7517), .B0(n1528), .B1(n7645), .Y(n5924) );
  OAI22XL U1290 ( .A0(n4139), .A1(n8029), .B0(n4150), .B1(n8157), .Y(n5922) );
  OAI22XL U1291 ( .A0(n4119), .A1(n7773), .B0(n4130), .B1(n7901), .Y(n5921) );
  OAI22XL U1292 ( .A0(n1704), .A1(n7518), .B0(n1528), .B1(n7646), .Y(n5928) );
  OAI22XL U1293 ( .A0(n4139), .A1(n8030), .B0(n4150), .B1(n8158), .Y(n5926) );
  OAI22XL U1294 ( .A0(n4119), .A1(n7774), .B0(n4130), .B1(n7902), .Y(n5925) );
  NOR4X1 U1295 ( .A(n1349), .B(n8274), .C(n6368), .D(n6367), .Y(n6369) );
  XOR2X1 U1296 ( .A(\tag_r[1][4] ), .B(n1312), .Y(n6368) );
  XOR2X1 U1297 ( .A(\tag_r[1][6] ), .B(n1314), .Y(n6367) );
  NOR4X1 U1298 ( .A(n3998), .B(n8273), .C(n6401), .D(n6400), .Y(n6402) );
  XOR2X1 U1299 ( .A(\tag_r[0][4] ), .B(n1312), .Y(n6401) );
  XOR2X1 U1300 ( .A(\tag_r[0][6] ), .B(n1314), .Y(n6400) );
  NOR4X1 U1301 ( .A(n1697), .B(n8275), .C(n6335), .D(n6334), .Y(n6336) );
  XOR2X1 U1302 ( .A(\tag_r[2][4] ), .B(n1312), .Y(n6335) );
  XOR2X1 U1303 ( .A(\tag_r[2][6] ), .B(n1314), .Y(n6334) );
  NOR4X1 U1304 ( .A(n1354), .B(n8276), .C(n6302), .D(n6301), .Y(n6303) );
  XOR2X1 U1305 ( .A(\tag_r[3][4] ), .B(n1312), .Y(n6302) );
  XOR2X1 U1306 ( .A(\tag_r[3][6] ), .B(n1314), .Y(n6301) );
  NAND4X1 U1307 ( .A(n6372), .B(n6371), .C(n6370), .D(n6369), .Y(n6399) );
  XOR2X1 U1308 ( .A(n7083), .B(n1319), .Y(n6372) );
  XOR2X1 U1309 ( .A(n7077), .B(n1313), .Y(n6371) );
  XOR2X1 U1310 ( .A(n7082), .B(n1318), .Y(n6370) );
  NAND4X1 U1311 ( .A(n6405), .B(n6404), .C(n6403), .D(n6402), .Y(n6432) );
  XOR2X1 U1312 ( .A(n7057), .B(n1318), .Y(n6405) );
  XOR2X1 U1313 ( .A(n7052), .B(n1313), .Y(n6404) );
  XOR2X1 U1314 ( .A(n7063), .B(n1324), .Y(n6403) );
  NAND4X1 U1315 ( .A(n6339), .B(n6338), .C(n6337), .D(n6336), .Y(n6366) );
  XOR2X1 U1316 ( .A(n7108), .B(n1319), .Y(n6339) );
  XOR2X1 U1317 ( .A(n7102), .B(n1313), .Y(n6338) );
  XOR2X1 U1318 ( .A(n7107), .B(n1318), .Y(n6337) );
  NAND4X1 U1319 ( .A(n6306), .B(n6305), .C(n6304), .D(n6303), .Y(n6333) );
  XOR2X1 U1320 ( .A(n7133), .B(n1319), .Y(n6306) );
  XOR2X1 U1321 ( .A(n7127), .B(n1313), .Y(n6305) );
  XOR2X1 U1322 ( .A(n7132), .B(n1318), .Y(n6304) );
  NAND3X1 U1323 ( .A(n6839), .B(n8271), .C(n6838), .Y(n7046) );
  NOR4X1 U1324 ( .A(n5757), .B(n5756), .C(n5755), .D(n5754), .Y(n5758) );
  OAI22XL U1325 ( .A0(n4134), .A1(n7197), .B0(n4149), .B1(n7222), .Y(n5757) );
  OAI22XL U1326 ( .A0(n4115), .A1(n7147), .B0(n4128), .B1(n7172), .Y(n5756) );
  NOR4X1 U1327 ( .A(n5762), .B(n5761), .C(n5760), .D(n5759), .Y(n5763) );
  OAI22XL U1328 ( .A0(n4134), .A1(n7198), .B0(n4149), .B1(n7223), .Y(n5762) );
  OAI22XL U1329 ( .A0(n4115), .A1(n7148), .B0(n4129), .B1(n7173), .Y(n5761) );
  NOR4X1 U1330 ( .A(n5767), .B(n5766), .C(n5765), .D(n5764), .Y(n5768) );
  OAI22XL U1331 ( .A0(n4134), .A1(n7199), .B0(n4149), .B1(n7224), .Y(n5767) );
  OAI22XL U1332 ( .A0(n4119), .A1(n7149), .B0(n4129), .B1(n7174), .Y(n5766) );
  NOR4X1 U1333 ( .A(n5772), .B(n5771), .C(n5770), .D(n5769), .Y(n5773) );
  OAI22XL U1334 ( .A0(n4134), .A1(n7200), .B0(n4149), .B1(n7225), .Y(n5772) );
  OAI22XL U1335 ( .A0(n4114), .A1(n7150), .B0(n4127), .B1(n7175), .Y(n5771) );
  NOR4X1 U1336 ( .A(n5777), .B(n5776), .C(n5775), .D(n5774), .Y(n5778) );
  OAI22XL U1337 ( .A0(n4141), .A1(n7201), .B0(n4151), .B1(n7226), .Y(n5777) );
  OAI22XL U1338 ( .A0(n4121), .A1(n7151), .B0(n4131), .B1(n7176), .Y(n5776) );
  NOR4X1 U1339 ( .A(n5782), .B(n5781), .C(n5780), .D(n5779), .Y(n5783) );
  OAI22XL U1340 ( .A0(n4141), .A1(n7202), .B0(n4151), .B1(n7227), .Y(n5782) );
  OAI22XL U1341 ( .A0(n4121), .A1(n7152), .B0(n4131), .B1(n7177), .Y(n5781) );
  NOR4X1 U1342 ( .A(n5787), .B(n5786), .C(n5785), .D(n5784), .Y(n5788) );
  OAI22XL U1343 ( .A0(n4141), .A1(n7203), .B0(n4151), .B1(n7228), .Y(n5787) );
  NOR4X1 U1344 ( .A(n5667), .B(n5666), .C(n5665), .D(n5664), .Y(n5668) );
  OAI22XL U1345 ( .A0(n4135), .A1(n7204), .B0(n4145), .B1(n7229), .Y(n5667) );
  OAI22XL U1346 ( .A0(n4115), .A1(n7154), .B0(n4125), .B1(n7179), .Y(n5666) );
  NOR4X1 U1347 ( .A(n5672), .B(n5671), .C(n5670), .D(n5669), .Y(n5673) );
  OAI22XL U1348 ( .A0(n4139), .A1(n7205), .B0(n4151), .B1(n7230), .Y(n5672) );
  OAI22XL U1349 ( .A0(n4121), .A1(n7155), .B0(n4127), .B1(n7180), .Y(n5671) );
  NOR4X1 U1350 ( .A(n5677), .B(n5676), .C(n5675), .D(n5674), .Y(n5678) );
  OAI22XL U1351 ( .A0(n4136), .A1(n7206), .B0(n4147), .B1(n7231), .Y(n5677) );
  OAI22XL U1352 ( .A0(n4114), .A1(n7156), .B0(n4131), .B1(n7181), .Y(n5676) );
  NOR4X1 U1353 ( .A(n5682), .B(n5681), .C(n5680), .D(n5679), .Y(n5683) );
  OAI22XL U1354 ( .A0(n4141), .A1(n7207), .B0(n4151), .B1(n7232), .Y(n5682) );
  OAI22XL U1355 ( .A0(n4121), .A1(n7157), .B0(n4127), .B1(n7182), .Y(n5681) );
  NOR4X1 U1356 ( .A(n5687), .B(n5686), .C(n5685), .D(n5684), .Y(n5688) );
  OAI22XL U1357 ( .A0(n4139), .A1(n7208), .B0(n4147), .B1(n7233), .Y(n5687) );
  OAI22XL U1358 ( .A0(n4114), .A1(n7158), .B0(n4131), .B1(n7183), .Y(n5686) );
  NOR4X1 U1359 ( .A(n5692), .B(n5691), .C(n5690), .D(n5689), .Y(n5693) );
  OAI22XL U1360 ( .A0(n4135), .A1(n7209), .B0(n4147), .B1(n7234), .Y(n5692) );
  OAI22XL U1361 ( .A0(n4114), .A1(n7159), .B0(n4129), .B1(n7184), .Y(n5691) );
  NOR4X1 U1362 ( .A(n5697), .B(n5696), .C(n5695), .D(n5694), .Y(n5698) );
  OAI22XL U1363 ( .A0(n6847), .A1(n7210), .B0(n4144), .B1(n7235), .Y(n5697) );
  OAI22XL U1364 ( .A0(n4114), .A1(n7160), .B0(n4128), .B1(n7185), .Y(n5696) );
  NOR4X1 U1365 ( .A(n5702), .B(n5701), .C(n5700), .D(n5699), .Y(n5703) );
  OAI22XL U1366 ( .A0(n6847), .A1(n7211), .B0(n4144), .B1(n7236), .Y(n5702) );
  OAI22XL U1367 ( .A0(n4114), .A1(n7161), .B0(n4128), .B1(n7186), .Y(n5701) );
  NOR4X1 U1368 ( .A(n5707), .B(n5706), .C(n5705), .D(n5704), .Y(n5708) );
  OAI22XL U1369 ( .A0(n6847), .A1(n7212), .B0(n4144), .B1(n7237), .Y(n5707) );
  OAI22XL U1370 ( .A0(n6845), .A1(n7162), .B0(n4128), .B1(n7187), .Y(n5706) );
  NOR4X1 U1371 ( .A(n5712), .B(n5711), .C(n5710), .D(n5709), .Y(n5713) );
  OAI22XL U1372 ( .A0(n6847), .A1(n7213), .B0(n4144), .B1(n7238), .Y(n5712) );
  OAI22XL U1373 ( .A0(n6845), .A1(n7163), .B0(n4124), .B1(n7188), .Y(n5711) );
  NOR4X1 U1374 ( .A(n5717), .B(n5716), .C(n5715), .D(n5714), .Y(n5718) );
  OAI22XL U1375 ( .A0(n6847), .A1(n7214), .B0(n4146), .B1(n7239), .Y(n5717) );
  OAI22XL U1376 ( .A0(n6845), .A1(n7164), .B0(n4124), .B1(n7189), .Y(n5716) );
  NOR4X1 U1377 ( .A(n5722), .B(n5721), .C(n5720), .D(n5719), .Y(n5723) );
  OAI22XL U1378 ( .A0(n6847), .A1(n7215), .B0(n4146), .B1(n7240), .Y(n5722) );
  OAI22XL U1379 ( .A0(n6845), .A1(n7165), .B0(n4124), .B1(n7190), .Y(n5721) );
  NOR4X1 U1380 ( .A(n5727), .B(n5726), .C(n5725), .D(n5724), .Y(n5728) );
  OAI22XL U1381 ( .A0(n4134), .A1(n7216), .B0(n4146), .B1(n7241), .Y(n5727) );
  OAI22XL U1382 ( .A0(n6845), .A1(n7166), .B0(n4126), .B1(n7191), .Y(n5726) );
  NOR4X1 U1383 ( .A(n5732), .B(n5731), .C(n5730), .D(n5729), .Y(n5733) );
  OAI22XL U1384 ( .A0(n4134), .A1(n7217), .B0(n4146), .B1(n7242), .Y(n5732) );
  OAI22XL U1385 ( .A0(n6845), .A1(n7167), .B0(n4126), .B1(n7192), .Y(n5731) );
  NOR4X1 U1386 ( .A(n5737), .B(n5736), .C(n5735), .D(n5734), .Y(n5738) );
  OAI22XL U1387 ( .A0(n4134), .A1(n7218), .B0(n4148), .B1(n7243), .Y(n5737) );
  OAI22XL U1388 ( .A0(n4114), .A1(n7168), .B0(n4124), .B1(n7193), .Y(n5736) );
  NOR4X1 U1389 ( .A(n5742), .B(n5741), .C(n5740), .D(n5739), .Y(n5743) );
  OAI22XL U1390 ( .A0(n4134), .A1(n7219), .B0(n4148), .B1(n7244), .Y(n5742) );
  OAI22XL U1391 ( .A0(n4114), .A1(n7169), .B0(n4129), .B1(n7194), .Y(n5741) );
  NOR4X1 U1392 ( .A(n5747), .B(n5746), .C(n5745), .D(n5744), .Y(n5748) );
  OAI22XL U1393 ( .A0(n4134), .A1(n7220), .B0(n4148), .B1(n7245), .Y(n5747) );
  OAI22XL U1394 ( .A0(n4114), .A1(n7170), .B0(n4126), .B1(n7195), .Y(n5746) );
  NOR4X1 U1395 ( .A(n5752), .B(n5751), .C(n5750), .D(n5749), .Y(n5753) );
  OAI22XL U1396 ( .A0(n4134), .A1(n7221), .B0(n4148), .B1(n7246), .Y(n5752) );
  OAI22XL U1397 ( .A0(n4114), .A1(n7171), .B0(n4126), .B1(n7196), .Y(n5751) );
  OAI22XL U1398 ( .A0(n4136), .A1(n8074), .B0(n4147), .B1(n8202), .Y(n6118) );
  OAI22XL U1399 ( .A0(n4116), .A1(n7818), .B0(n4127), .B1(n7946), .Y(n6117) );
  OAI22XL U1400 ( .A0(n1701), .A1(n7562), .B0(n1358), .B1(n7690), .Y(n6120) );
  OAI22XL U1401 ( .A0(n4136), .A1(n8075), .B0(n4147), .B1(n8203), .Y(n6126) );
  OAI22XL U1402 ( .A0(n4116), .A1(n7819), .B0(n4127), .B1(n7947), .Y(n6125) );
  OAI22XL U1403 ( .A0(n1701), .A1(n7563), .B0(n1358), .B1(n7691), .Y(n6128) );
  OAI22XL U1404 ( .A0(n4138), .A1(n8094), .B0(n4146), .B1(n8222), .Y(n6206) );
  OAI22XL U1405 ( .A0(n4118), .A1(n7838), .B0(n4126), .B1(n7966), .Y(n6205) );
  OAI22XL U1406 ( .A0(n1695), .A1(n7582), .B0(n1357), .B1(n7710), .Y(n6208) );
  OAI22XL U1407 ( .A0(n4135), .A1(n8106), .B0(n4145), .B1(n8234), .Y(n6262) );
  OAI22XL U1408 ( .A0(n4115), .A1(n7850), .B0(n4125), .B1(n7978), .Y(n6261) );
  OAI22XL U1409 ( .A0(n1697), .A1(n7594), .B0(n1355), .B1(n7722), .Y(n6264) );
  OAI22XL U1410 ( .A0(n4135), .A1(n8107), .B0(n4145), .B1(n8235), .Y(n6266) );
  OAI22XL U1411 ( .A0(n4115), .A1(n7851), .B0(n4125), .B1(n7979), .Y(n6265) );
  OAI22XL U1412 ( .A0(n1697), .A1(n7595), .B0(n1359), .B1(n7723), .Y(n6268) );
  OAI22XL U1413 ( .A0(n4140), .A1(n8138), .B0(n4145), .B1(n8266), .Y(n5894) );
  OAI22XL U1414 ( .A0(n4120), .A1(n7882), .B0(n4125), .B1(n8010), .Y(n5893) );
  OAI22XL U1415 ( .A0(n1696), .A1(n7626), .B0(n1580), .B1(n7754), .Y(n5896) );
  OAI22XL U1416 ( .A0(n4140), .A1(n8139), .B0(n4150), .B1(n8267), .Y(n5898) );
  OAI22XL U1417 ( .A0(n4120), .A1(n7883), .B0(n4130), .B1(n8011), .Y(n5897) );
  OAI22XL U1418 ( .A0(n1703), .A1(n7627), .B0(n1356), .B1(n7755), .Y(n5900) );
  OAI22XL U1419 ( .A0(n4139), .A1(n8042), .B0(n4150), .B1(n8170), .Y(n5978) );
  OAI22XL U1420 ( .A0(n4119), .A1(n7786), .B0(n4130), .B1(n7914), .Y(n5977) );
  OAI22XL U1421 ( .A0(n1704), .A1(n7530), .B0(n1528), .B1(n7658), .Y(n5980) );
  OAI22XL U1422 ( .A0(n4138), .A1(n8043), .B0(n4149), .B1(n8171), .Y(n5982) );
  OAI22XL U1423 ( .A0(n4118), .A1(n7787), .B0(n4129), .B1(n7915), .Y(n5981) );
  OAI22XL U1424 ( .A0(n1703), .A1(n7531), .B0(n1359), .B1(n7659), .Y(n5984) );
  XOR2X1 U1425 ( .A(\tag_r[1][3] ), .B(n1311), .Y(n6381) );
  XOR2X1 U1426 ( .A(\tag_r[1][17] ), .B(n1325), .Y(n6373) );
  XOR2X1 U1427 ( .A(\tag_r[0][3] ), .B(n1311), .Y(n6414) );
  XOR2X1 U1428 ( .A(\tag_r[0][17] ), .B(n1325), .Y(n6406) );
  XOR2X1 U1429 ( .A(\tag_r[2][3] ), .B(n1311), .Y(n6348) );
  XOR2X1 U1430 ( .A(\tag_r[2][17] ), .B(n1325), .Y(n6340) );
  XOR2X1 U1431 ( .A(\tag_r[3][3] ), .B(n1311), .Y(n6315) );
  XOR2X1 U1432 ( .A(\tag_r[3][17] ), .B(n1325), .Y(n6307) );
  XOR2X1 U1433 ( .A(\tag_r[5][3] ), .B(n1311), .Y(n6517) );
  XOR2X1 U1434 ( .A(\tag_r[5][17] ), .B(n1325), .Y(n6509) );
  XOR2X1 U1435 ( .A(\tag_r[4][3] ), .B(n1311), .Y(n6550) );
  XOR2X1 U1436 ( .A(\tag_r[4][17] ), .B(n1325), .Y(n6542) );
  XOR2X1 U1437 ( .A(\tag_r[6][3] ), .B(n1311), .Y(n6484) );
  XOR2X1 U1438 ( .A(\tag_r[6][17] ), .B(n1325), .Y(n6476) );
  XOR2X1 U1439 ( .A(\tag_r[7][3] ), .B(n1311), .Y(n6451) );
  XOR2X1 U1440 ( .A(\tag_r[7][17] ), .B(n1325), .Y(n6443) );
  NOR4X1 U1441 ( .A(n6384), .B(n6383), .C(n6382), .D(n6381), .Y(n6385) );
  XOR2X1 U1442 ( .A(\tag_r[1][0] ), .B(n1308), .Y(n6384) );
  XOR2X1 U1443 ( .A(\tag_r[1][1] ), .B(n1309), .Y(n6383) );
  XOR2X1 U1444 ( .A(\tag_r[1][2] ), .B(n1310), .Y(n6382) );
  NOR4X1 U1445 ( .A(n6376), .B(n6375), .C(n6374), .D(n6373), .Y(n6377) );
  XOR2X1 U1446 ( .A(\tag_r[1][12] ), .B(n1320), .Y(n6376) );
  XOR2X1 U1447 ( .A(\tag_r[1][16] ), .B(n1324), .Y(n6375) );
  XOR2X1 U1448 ( .A(\tag_r[1][18] ), .B(n1326), .Y(n6374) );
  NOR4X1 U1449 ( .A(n6417), .B(n6416), .C(n6415), .D(n6414), .Y(n6418) );
  XOR2X1 U1450 ( .A(\tag_r[0][0] ), .B(n1308), .Y(n6417) );
  XOR2X1 U1451 ( .A(\tag_r[0][1] ), .B(n1309), .Y(n6416) );
  XOR2X1 U1452 ( .A(\tag_r[0][2] ), .B(n1310), .Y(n6415) );
  NOR4X1 U1453 ( .A(n6409), .B(n6408), .C(n6407), .D(n6406), .Y(n6410) );
  XOR2X1 U1454 ( .A(\tag_r[0][12] ), .B(n1320), .Y(n6409) );
  XOR2X1 U1455 ( .A(\tag_r[0][11] ), .B(n1319), .Y(n6408) );
  XOR2X1 U1456 ( .A(\tag_r[0][18] ), .B(n1326), .Y(n6407) );
  NOR4X1 U1457 ( .A(n6351), .B(n6350), .C(n6349), .D(n6348), .Y(n6352) );
  XOR2X1 U1458 ( .A(\tag_r[2][0] ), .B(n1308), .Y(n6351) );
  XOR2X1 U1459 ( .A(\tag_r[2][1] ), .B(n1309), .Y(n6350) );
  XOR2X1 U1460 ( .A(\tag_r[2][2] ), .B(n1310), .Y(n6349) );
  NOR4X1 U1461 ( .A(n6343), .B(n6342), .C(n6341), .D(n6340), .Y(n6344) );
  XOR2X1 U1462 ( .A(\tag_r[2][12] ), .B(n1320), .Y(n6343) );
  XOR2X1 U1463 ( .A(\tag_r[2][16] ), .B(n1324), .Y(n6342) );
  XOR2X1 U1464 ( .A(\tag_r[2][18] ), .B(n1326), .Y(n6341) );
  NOR4X1 U1465 ( .A(n6318), .B(n6317), .C(n6316), .D(n6315), .Y(n6319) );
  XOR2X1 U1466 ( .A(\tag_r[3][0] ), .B(n1308), .Y(n6318) );
  XOR2X1 U1467 ( .A(\tag_r[3][1] ), .B(n1309), .Y(n6317) );
  XOR2X1 U1468 ( .A(\tag_r[3][2] ), .B(n1310), .Y(n6316) );
  NOR4X1 U1469 ( .A(n6310), .B(n6309), .C(n6308), .D(n6307), .Y(n6311) );
  XOR2X1 U1470 ( .A(\tag_r[3][12] ), .B(n1320), .Y(n6310) );
  XOR2X1 U1471 ( .A(\tag_r[3][16] ), .B(n1324), .Y(n6309) );
  XOR2X1 U1472 ( .A(\tag_r[3][18] ), .B(n1326), .Y(n6308) );
  NOR4X1 U1473 ( .A(n4125), .B(n8278), .C(n6504), .D(n6503), .Y(n6505) );
  XOR2X1 U1474 ( .A(\tag_r[5][4] ), .B(n1312), .Y(n6504) );
  XOR2X1 U1475 ( .A(\tag_r[5][6] ), .B(n1314), .Y(n6503) );
  NOR4X1 U1476 ( .A(n6520), .B(n6519), .C(n6518), .D(n6517), .Y(n6521) );
  XOR2X1 U1477 ( .A(\tag_r[5][0] ), .B(n1308), .Y(n6520) );
  XOR2X1 U1478 ( .A(\tag_r[5][1] ), .B(n1309), .Y(n6519) );
  XOR2X1 U1479 ( .A(\tag_r[5][2] ), .B(n1310), .Y(n6518) );
  NOR4X1 U1480 ( .A(n6512), .B(n6511), .C(n6510), .D(n6509), .Y(n6513) );
  XOR2X1 U1481 ( .A(\tag_r[5][12] ), .B(n1320), .Y(n6512) );
  XOR2X1 U1482 ( .A(\tag_r[5][16] ), .B(n1324), .Y(n6511) );
  XOR2X1 U1483 ( .A(\tag_r[5][18] ), .B(n1326), .Y(n6510) );
  NOR4X1 U1484 ( .A(n4115), .B(n8277), .C(n6537), .D(n6536), .Y(n6538) );
  XOR2X1 U1485 ( .A(\tag_r[4][4] ), .B(n1312), .Y(n6537) );
  XOR2X1 U1486 ( .A(\tag_r[4][6] ), .B(n1314), .Y(n6536) );
  NOR4X1 U1487 ( .A(n6553), .B(n6552), .C(n6551), .D(n6550), .Y(n6554) );
  XOR2X1 U1488 ( .A(\tag_r[4][0] ), .B(n1308), .Y(n6553) );
  XOR2X1 U1489 ( .A(\tag_r[4][1] ), .B(n1309), .Y(n6552) );
  XOR2X1 U1490 ( .A(\tag_r[4][2] ), .B(n1310), .Y(n6551) );
  NOR4X1 U1491 ( .A(n6545), .B(n6544), .C(n6543), .D(n6542), .Y(n6546) );
  XOR2X1 U1492 ( .A(\tag_r[4][12] ), .B(n1320), .Y(n6545) );
  XOR2X1 U1493 ( .A(\tag_r[4][16] ), .B(n1324), .Y(n6544) );
  XOR2X1 U1494 ( .A(\tag_r[4][18] ), .B(n1326), .Y(n6543) );
  NOR4X1 U1495 ( .A(n4135), .B(n8279), .C(n6471), .D(n6470), .Y(n6472) );
  XOR2X1 U1496 ( .A(\tag_r[6][4] ), .B(n1312), .Y(n6471) );
  XOR2X1 U1497 ( .A(\tag_r[6][6] ), .B(n1314), .Y(n6470) );
  NOR4X1 U1498 ( .A(n6487), .B(n6486), .C(n6485), .D(n6484), .Y(n6488) );
  XOR2X1 U1499 ( .A(\tag_r[6][0] ), .B(n1308), .Y(n6487) );
  XOR2X1 U1500 ( .A(\tag_r[6][1] ), .B(n1309), .Y(n6486) );
  XOR2X1 U1501 ( .A(\tag_r[6][2] ), .B(n1310), .Y(n6485) );
  NOR4X1 U1502 ( .A(n6479), .B(n6478), .C(n6477), .D(n6476), .Y(n6480) );
  XOR2X1 U1503 ( .A(\tag_r[6][12] ), .B(n1320), .Y(n6479) );
  XOR2X1 U1504 ( .A(\tag_r[6][16] ), .B(n1324), .Y(n6478) );
  XOR2X1 U1505 ( .A(\tag_r[6][18] ), .B(n1326), .Y(n6477) );
  NOR4X1 U1506 ( .A(n4145), .B(n8280), .C(n6438), .D(n6437), .Y(n6439) );
  XOR2X1 U1507 ( .A(\tag_r[7][4] ), .B(n1312), .Y(n6438) );
  XOR2X1 U1508 ( .A(\tag_r[7][6] ), .B(n1314), .Y(n6437) );
  NOR4X1 U1509 ( .A(n6454), .B(n6453), .C(n6452), .D(n6451), .Y(n6455) );
  XOR2X1 U1510 ( .A(\tag_r[7][0] ), .B(n1308), .Y(n6454) );
  XOR2X1 U1511 ( .A(\tag_r[7][1] ), .B(n1309), .Y(n6453) );
  XOR2X1 U1512 ( .A(\tag_r[7][2] ), .B(n1310), .Y(n6452) );
  NOR4X1 U1513 ( .A(n6446), .B(n6445), .C(n6444), .D(n6443), .Y(n6447) );
  XOR2X1 U1514 ( .A(\tag_r[7][12] ), .B(n1320), .Y(n6446) );
  XOR2X1 U1515 ( .A(\tag_r[7][11] ), .B(n1319), .Y(n6445) );
  XOR2X1 U1516 ( .A(\tag_r[7][18] ), .B(n1326), .Y(n6444) );
  XOR2X1 U1517 ( .A(n7081), .B(n1317), .Y(n6386) );
  XOR2X1 U1518 ( .A(n7095), .B(n1331), .Y(n6378) );
  XOR2X1 U1519 ( .A(n7093), .B(n1329), .Y(n6393) );
  XOR2X1 U1520 ( .A(n7056), .B(n1317), .Y(n6419) );
  XOR2X1 U1521 ( .A(n7070), .B(n1331), .Y(n6411) );
  XOR2X1 U1522 ( .A(n7068), .B(n1329), .Y(n6426) );
  XOR2X1 U1523 ( .A(n7106), .B(n1317), .Y(n6353) );
  XOR2X1 U1524 ( .A(n7120), .B(n1331), .Y(n6345) );
  XOR2X1 U1525 ( .A(n7118), .B(n1329), .Y(n6360) );
  XOR2X1 U1526 ( .A(n7131), .B(n1317), .Y(n6320) );
  XOR2X1 U1527 ( .A(n7145), .B(n1331), .Y(n6312) );
  XOR2X1 U1528 ( .A(n7143), .B(n1329), .Y(n6327) );
  XOR2X1 U1529 ( .A(n7181), .B(n1317), .Y(n6522) );
  XOR2X1 U1530 ( .A(n7195), .B(n1331), .Y(n6514) );
  XOR2X1 U1531 ( .A(n7193), .B(n1329), .Y(n6529) );
  XOR2X1 U1532 ( .A(n7156), .B(n1317), .Y(n6555) );
  XOR2X1 U1533 ( .A(n7170), .B(n1331), .Y(n6547) );
  XOR2X1 U1534 ( .A(n7168), .B(n1329), .Y(n6562) );
  XOR2X1 U1535 ( .A(n7206), .B(n1317), .Y(n6489) );
  XOR2X1 U1536 ( .A(n7220), .B(n1331), .Y(n6481) );
  XOR2X1 U1537 ( .A(n7218), .B(n1329), .Y(n6496) );
  XOR2X1 U1538 ( .A(n7079), .B(n1315), .Y(n6387) );
  XOR2X1 U1539 ( .A(n7094), .B(n1330), .Y(n6379) );
  XOR2X1 U1540 ( .A(n7091), .B(n1327), .Y(n6394) );
  XOR2X1 U1541 ( .A(n7054), .B(n1315), .Y(n6420) );
  XOR2X1 U1542 ( .A(n7069), .B(n1330), .Y(n6412) );
  XOR2X1 U1543 ( .A(n7066), .B(n1327), .Y(n6427) );
  XOR2X1 U1544 ( .A(n7104), .B(n1315), .Y(n6354) );
  XOR2X1 U1545 ( .A(n7119), .B(n1330), .Y(n6346) );
  XOR2X1 U1546 ( .A(n7116), .B(n1327), .Y(n6361) );
  XOR2X1 U1547 ( .A(n7129), .B(n1315), .Y(n6321) );
  XOR2X1 U1548 ( .A(n7144), .B(n1330), .Y(n6313) );
  XOR2X1 U1549 ( .A(n7141), .B(n1327), .Y(n6328) );
  XOR2X1 U1550 ( .A(n7179), .B(n1315), .Y(n6523) );
  XOR2X1 U1551 ( .A(n7194), .B(n1330), .Y(n6515) );
  XOR2X1 U1552 ( .A(n7191), .B(n1327), .Y(n6530) );
  XOR2X1 U1553 ( .A(n7154), .B(n1315), .Y(n6556) );
  XOR2X1 U1554 ( .A(n7169), .B(n1330), .Y(n6548) );
  XOR2X1 U1555 ( .A(n7166), .B(n1327), .Y(n6563) );
  XOR2X1 U1556 ( .A(n7204), .B(n1315), .Y(n6490) );
  XOR2X1 U1557 ( .A(n7219), .B(n1330), .Y(n6482) );
  XOR2X1 U1558 ( .A(n7216), .B(n1327), .Y(n6497) );
  XOR2X1 U1559 ( .A(n7080), .B(n1316), .Y(n6388) );
  XOR2X1 U1560 ( .A(n7096), .B(n1332), .Y(n6380) );
  XOR2X1 U1561 ( .A(n7092), .B(n1328), .Y(n6395) );
  XOR2X1 U1562 ( .A(n7055), .B(n1316), .Y(n6421) );
  XOR2X1 U1563 ( .A(n7071), .B(n1332), .Y(n6413) );
  XOR2X1 U1564 ( .A(n7067), .B(n1328), .Y(n6428) );
  XOR2X1 U1565 ( .A(n7105), .B(n1316), .Y(n6355) );
  XOR2X1 U1566 ( .A(n7121), .B(n1332), .Y(n6347) );
  XOR2X1 U1567 ( .A(n7117), .B(n1328), .Y(n6362) );
  XOR2X1 U1568 ( .A(n7130), .B(n1316), .Y(n6322) );
  XOR2X1 U1569 ( .A(n7146), .B(n1332), .Y(n6314) );
  XOR2X1 U1570 ( .A(n7142), .B(n1328), .Y(n6329) );
  XOR2X1 U1571 ( .A(n7180), .B(n1316), .Y(n6524) );
  XOR2X1 U1572 ( .A(n7196), .B(n1332), .Y(n6516) );
  XOR2X1 U1573 ( .A(n7192), .B(n1328), .Y(n6531) );
  XOR2X1 U1574 ( .A(n7155), .B(n1316), .Y(n6557) );
  XOR2X1 U1575 ( .A(n7171), .B(n1332), .Y(n6549) );
  XOR2X1 U1576 ( .A(n7167), .B(n1328), .Y(n6564) );
  XOR2X1 U1577 ( .A(n7205), .B(n1316), .Y(n6491) );
  XOR2X1 U1578 ( .A(n7221), .B(n1332), .Y(n6483) );
  XOR2X1 U1579 ( .A(n7217), .B(n1328), .Y(n6498) );
  NAND4X1 U1580 ( .A(n6465), .B(n6464), .C(n6463), .D(n6462), .Y(n6466) );
  XOR2X1 U1581 ( .A(n7242), .B(n1328), .Y(n6465) );
  XOR2X1 U1582 ( .A(n7241), .B(n1327), .Y(n6464) );
  XOR2X1 U1583 ( .A(n7243), .B(n1329), .Y(n6463) );
  NAND4X1 U1584 ( .A(n6458), .B(n6457), .C(n6456), .D(n6455), .Y(n6467) );
  XOR2X1 U1585 ( .A(n7230), .B(n1316), .Y(n6458) );
  XOR2X1 U1586 ( .A(n7229), .B(n1315), .Y(n6457) );
  XOR2X1 U1587 ( .A(n7231), .B(n1317), .Y(n6456) );
  NAND4X1 U1588 ( .A(n6508), .B(n6507), .C(n6506), .D(n6505), .Y(n6535) );
  XOR2X1 U1589 ( .A(n7183), .B(n1319), .Y(n6508) );
  XOR2X1 U1590 ( .A(n7177), .B(n1313), .Y(n6507) );
  XOR2X1 U1591 ( .A(n7182), .B(n1318), .Y(n6506) );
  NAND4X1 U1592 ( .A(n6541), .B(n6540), .C(n6539), .D(n6538), .Y(n6568) );
  XOR2X1 U1593 ( .A(n7158), .B(n1319), .Y(n6541) );
  XOR2X1 U1594 ( .A(n7152), .B(n1313), .Y(n6540) );
  XOR2X1 U1595 ( .A(n7157), .B(n1318), .Y(n6539) );
  NAND4X1 U1596 ( .A(n6475), .B(n6474), .C(n6473), .D(n6472), .Y(n6502) );
  XOR2X1 U1597 ( .A(n7208), .B(n1319), .Y(n6475) );
  XOR2X1 U1598 ( .A(n7202), .B(n1313), .Y(n6474) );
  XOR2X1 U1599 ( .A(n7207), .B(n1318), .Y(n6473) );
  NAND4X1 U1600 ( .A(n6442), .B(n6441), .C(n6440), .D(n6439), .Y(n6469) );
  XOR2X1 U1601 ( .A(n7232), .B(n1318), .Y(n6442) );
  XOR2X1 U1602 ( .A(n7227), .B(n1313), .Y(n6441) );
  XOR2X1 U1603 ( .A(n7238), .B(n1324), .Y(n6440) );
  NAND4X1 U1604 ( .A(n6450), .B(n6449), .C(n6448), .D(n6447), .Y(n6468) );
  XOR2X1 U1605 ( .A(n7246), .B(n1332), .Y(n6450) );
  XOR2X1 U1606 ( .A(n7244), .B(n1330), .Y(n6449) );
  XOR2X1 U1607 ( .A(n7245), .B(n1331), .Y(n6448) );
  NOR3X1 U1608 ( .A(n6391), .B(n6390), .C(n6389), .Y(n6392) );
  XOR2X1 U1609 ( .A(\tag_r[1][15] ), .B(n1323), .Y(n6391) );
  XOR2X1 U1610 ( .A(\tag_r[1][13] ), .B(n1321), .Y(n6390) );
  XOR2X1 U1611 ( .A(\tag_r[1][14] ), .B(n1322), .Y(n6389) );
  NOR3X1 U1612 ( .A(n6424), .B(n6423), .C(n6422), .Y(n6425) );
  XOR2X1 U1613 ( .A(\tag_r[0][15] ), .B(n1323), .Y(n6424) );
  XOR2X1 U1614 ( .A(\tag_r[0][13] ), .B(n1321), .Y(n6423) );
  XOR2X1 U1615 ( .A(\tag_r[0][14] ), .B(n1322), .Y(n6422) );
  NOR3X1 U1616 ( .A(n6358), .B(n6357), .C(n6356), .Y(n6359) );
  XOR2X1 U1617 ( .A(\tag_r[2][15] ), .B(n1323), .Y(n6358) );
  XOR2X1 U1618 ( .A(\tag_r[2][13] ), .B(n1321), .Y(n6357) );
  XOR2X1 U1619 ( .A(\tag_r[2][14] ), .B(n1322), .Y(n6356) );
  NOR3X1 U1620 ( .A(n6325), .B(n6324), .C(n6323), .Y(n6326) );
  XOR2X1 U1621 ( .A(\tag_r[3][15] ), .B(n1323), .Y(n6325) );
  XOR2X1 U1622 ( .A(\tag_r[3][13] ), .B(n1321), .Y(n6324) );
  XOR2X1 U1623 ( .A(\tag_r[3][14] ), .B(n1322), .Y(n6323) );
  NOR3X1 U1624 ( .A(n6527), .B(n6526), .C(n6525), .Y(n6528) );
  XOR2X1 U1625 ( .A(\tag_r[5][15] ), .B(n1323), .Y(n6527) );
  XOR2X1 U1626 ( .A(\tag_r[5][13] ), .B(n1321), .Y(n6526) );
  XOR2X1 U1627 ( .A(\tag_r[5][14] ), .B(n1322), .Y(n6525) );
  NOR3X1 U1628 ( .A(n6560), .B(n6559), .C(n6558), .Y(n6561) );
  XOR2X1 U1629 ( .A(\tag_r[4][15] ), .B(n1323), .Y(n6560) );
  XOR2X1 U1630 ( .A(\tag_r[4][13] ), .B(n1321), .Y(n6559) );
  XOR2X1 U1631 ( .A(\tag_r[4][14] ), .B(n1322), .Y(n6558) );
  NOR3X1 U1632 ( .A(n6494), .B(n6493), .C(n6492), .Y(n6495) );
  XOR2X1 U1633 ( .A(\tag_r[6][15] ), .B(n1323), .Y(n6494) );
  XOR2X1 U1634 ( .A(\tag_r[6][13] ), .B(n1321), .Y(n6493) );
  XOR2X1 U1635 ( .A(\tag_r[6][14] ), .B(n1322), .Y(n6492) );
  NOR3X1 U1636 ( .A(n6461), .B(n6460), .C(n6459), .Y(n6462) );
  XOR2X1 U1637 ( .A(\tag_r[7][15] ), .B(n1323), .Y(n6461) );
  XOR2X1 U1638 ( .A(\tag_r[7][13] ), .B(n1321), .Y(n6460) );
  XOR2X1 U1639 ( .A(\tag_r[7][14] ), .B(n1322), .Y(n6459) );
  CLKBUFX3 U1640 ( .A(proc_addr[11]), .Y(n1314) );
  CLKBUFX3 U1641 ( .A(proc_addr[9]), .Y(n1312) );
  CLKBUFX3 U1642 ( .A(proc_addr[8]), .Y(n1311) );
  CLKBUFX3 U1643 ( .A(proc_addr[7]), .Y(n1310) );
  CLKBUFX3 U1644 ( .A(proc_addr[6]), .Y(n1309) );
  CLKBUFX3 U1645 ( .A(proc_addr[5]), .Y(n1308) );
  CLKBUFX3 U1646 ( .A(proc_addr[22]), .Y(n1325) );
  CLKBUFX3 U1647 ( .A(proc_addr[23]), .Y(n1326) );
  CLKBUFX3 U1648 ( .A(proc_addr[17]), .Y(n1320) );
  CLKBUFX3 U1649 ( .A(proc_addr[19]), .Y(n1322) );
  CLKBUFX3 U1650 ( .A(proc_addr[18]), .Y(n1321) );
  CLKBUFX3 U1651 ( .A(proc_addr[20]), .Y(n1323) );
  CLKBUFX3 U1652 ( .A(proc_addr[16]), .Y(n1319) );
  CLKBUFX3 U1653 ( .A(proc_addr[21]), .Y(n1324) );
  CLKBUFX3 U1654 ( .A(proc_addr[10]), .Y(n1313) );
  CLKBUFX3 U1655 ( .A(proc_addr[15]), .Y(n1318) );
  CLKBUFX3 U1656 ( .A(proc_addr[14]), .Y(n1317) );
  CLKBUFX3 U1657 ( .A(proc_addr[12]), .Y(n1315) );
  CLKBUFX3 U1658 ( .A(proc_addr[13]), .Y(n1316) );
  CLKBUFX3 U1659 ( .A(proc_addr[28]), .Y(n1331) );
  CLKBUFX3 U1660 ( .A(proc_addr[27]), .Y(n1330) );
  CLKBUFX3 U1661 ( .A(proc_addr[26]), .Y(n1329) );
  CLKBUFX3 U1662 ( .A(proc_addr[24]), .Y(n1327) );
  CLKBUFX3 U1663 ( .A(proc_addr[25]), .Y(n1328) );
  CLKBUFX3 U1664 ( .A(proc_addr[29]), .Y(n1332) );
  AOI22X2 U1665 ( .A0(mem_rdata[19]), .A1(n1345), .B0(n4010), .B1(n6576), .Y(
        n6720) );
  OAI22XL U1666 ( .A0(n4196), .A1(n4375), .B0(n6932), .B1(n6706), .Y(n6576) );
  AOI22X2 U1667 ( .A0(mem_rdata[20]), .A1(n1345), .B0(n4010), .B1(n6577), .Y(
        n6721) );
  OAI22XL U1668 ( .A0(n4196), .A1(n4376), .B0(n6942), .B1(n6706), .Y(n6577) );
  AOI22X2 U1669 ( .A0(mem_rdata[21]), .A1(n1345), .B0(n4010), .B1(n6578), .Y(
        n6722) );
  OAI22XL U1670 ( .A0(n4196), .A1(n4377), .B0(n6947), .B1(n6706), .Y(n6578) );
  AOI22X2 U1671 ( .A0(mem_rdata[22]), .A1(n1345), .B0(n4010), .B1(n6579), .Y(
        n6723) );
  OAI22XL U1672 ( .A0(n4196), .A1(n4378), .B0(n6952), .B1(n6706), .Y(n6579) );
  AOI22X2 U1673 ( .A0(mem_rdata[23]), .A1(n1345), .B0(n4010), .B1(n6580), .Y(
        n6724) );
  OAI22XL U1674 ( .A0(n7038), .A1(n4379), .B0(n6957), .B1(n4009), .Y(n6580) );
  AOI22X2 U1675 ( .A0(mem_rdata[24]), .A1(n1345), .B0(n4010), .B1(n6581), .Y(
        n6725) );
  OAI22XL U1676 ( .A0(n4196), .A1(n4380), .B0(n6962), .B1(n4009), .Y(n6581) );
  AOI22X2 U1677 ( .A0(mem_rdata[25]), .A1(n1345), .B0(n4010), .B1(n6582), .Y(
        n6726) );
  OAI22XL U1678 ( .A0(n4196), .A1(n4381), .B0(n6967), .B1(n4009), .Y(n6582) );
  AOI22X2 U1679 ( .A0(mem_rdata[26]), .A1(n1345), .B0(n4010), .B1(n6583), .Y(
        n6727) );
  OAI22XL U1680 ( .A0(n4196), .A1(n4382), .B0(n6972), .B1(n4009), .Y(n6583) );
  AOI22X2 U1681 ( .A0(mem_rdata[27]), .A1(n4351), .B0(n4010), .B1(n6584), .Y(
        n6728) );
  OAI22XL U1682 ( .A0(n4196), .A1(n4383), .B0(n6977), .B1(n4009), .Y(n6584) );
  AOI22X2 U1683 ( .A0(mem_rdata[28]), .A1(n1338), .B0(n4010), .B1(n6585), .Y(
        n6729) );
  OAI22XL U1684 ( .A0(n7038), .A1(n4384), .B0(n6982), .B1(n4009), .Y(n6585) );
  AOI22X2 U1685 ( .A0(mem_rdata[29]), .A1(n1340), .B0(n4010), .B1(n6586), .Y(
        n6730) );
  OAI22XL U1686 ( .A0(n7038), .A1(n4385), .B0(n6987), .B1(n4009), .Y(n6586) );
  AOI22X2 U1687 ( .A0(mem_rdata[30]), .A1(n1341), .B0(n4011), .B1(n6587), .Y(
        n6731) );
  OAI22XL U1688 ( .A0(n4195), .A1(n4386), .B0(n6997), .B1(n4009), .Y(n6587) );
  AOI22X2 U1689 ( .A0(mem_rdata[31]), .A1(n1343), .B0(n4011), .B1(n6588), .Y(
        n6732) );
  OAI22XL U1690 ( .A0(n4195), .A1(n4387), .B0(n7002), .B1(n4009), .Y(n6588) );
  AOI22X2 U1691 ( .A0(mem_rdata[32]), .A1(n1342), .B0(n4011), .B1(n6589), .Y(
        n6733) );
  OAI22XL U1692 ( .A0(n4199), .A1(n4356), .B0(n6884), .B1(n4006), .Y(n6589) );
  AOI22X2 U1693 ( .A0(mem_rdata[33]), .A1(n1344), .B0(n4011), .B1(n6590), .Y(
        n6734) );
  OAI22XL U1694 ( .A0(n4200), .A1(n4357), .B0(n6939), .B1(n4006), .Y(n6590) );
  AOI22X2 U1695 ( .A0(mem_rdata[34]), .A1(n1339), .B0(n4011), .B1(n6591), .Y(
        n6735) );
  OAI22XL U1696 ( .A0(n4198), .A1(n4358), .B0(n6994), .B1(n4006), .Y(n6591) );
  AOI22X2 U1697 ( .A0(mem_rdata[89]), .A1(n1341), .B0(n4014), .B1(n6648), .Y(
        n6790) );
  OAI22XL U1698 ( .A0(n4203), .A1(n4381), .B0(n6970), .B1(n6654), .Y(n6648) );
  AOI22X2 U1699 ( .A0(mem_rdata[90]), .A1(n1341), .B0(n4015), .B1(n6649), .Y(
        n6791) );
  OAI22XL U1700 ( .A0(n4202), .A1(n4382), .B0(n6975), .B1(n6654), .Y(n6649) );
  AOI22X2 U1701 ( .A0(mem_rdata[91]), .A1(n1341), .B0(n4015), .B1(n6650), .Y(
        n6792) );
  OAI22XL U1702 ( .A0(n4203), .A1(n4383), .B0(n6980), .B1(n6654), .Y(n6650) );
  AOI22X2 U1703 ( .A0(mem_rdata[92]), .A1(n1341), .B0(n4015), .B1(n6651), .Y(
        n6793) );
  OAI22XL U1704 ( .A0(n4202), .A1(n4384), .B0(n6985), .B1(n6654), .Y(n6651) );
  AOI22X2 U1705 ( .A0(mem_rdata[93]), .A1(n1341), .B0(n4015), .B1(n6652), .Y(
        n6794) );
  OAI22XL U1706 ( .A0(n4205), .A1(n4385), .B0(n6990), .B1(n6654), .Y(n6652) );
  AOI22X2 U1707 ( .A0(mem_rdata[94]), .A1(n1341), .B0(n4015), .B1(n6653), .Y(
        n6795) );
  OAI22XL U1708 ( .A0(n4202), .A1(n4386), .B0(n7000), .B1(n6654), .Y(n6653) );
  AOI22X2 U1709 ( .A0(mem_rdata[95]), .A1(n1341), .B0(n4015), .B1(n6655), .Y(
        n6796) );
  OAI22XL U1710 ( .A0(n4202), .A1(n4387), .B0(n7005), .B1(n6654), .Y(n6655) );
  AOI22X2 U1711 ( .A0(mem_rdata[96]), .A1(n1341), .B0(n4015), .B1(n6656), .Y(
        n6797) );
  OAI22XL U1712 ( .A0(n6881), .A1(n6687), .B0(n4193), .B1(n4356), .Y(n6656) );
  AOI22X2 U1713 ( .A0(mem_rdata[97]), .A1(n1341), .B0(n4015), .B1(n6657), .Y(
        n6798) );
  OAI22XL U1714 ( .A0(n6936), .A1(n6687), .B0(n4193), .B1(n4357), .Y(n6657) );
  AOI22X2 U1715 ( .A0(mem_rdata[98]), .A1(n1340), .B0(n4015), .B1(n6658), .Y(
        n6799) );
  OAI22XL U1716 ( .A0(n6991), .A1(n4008), .B0(n4193), .B1(n4358), .Y(n6658) );
  AOI22X2 U1717 ( .A0(mem_rdata[99]), .A1(n1340), .B0(n4015), .B1(n6659), .Y(
        n6800) );
  OAI22XL U1718 ( .A0(n7006), .A1(n4008), .B0(n4193), .B1(n4359), .Y(n6659) );
  AOI22X2 U1719 ( .A0(mem_rdata[100]), .A1(n1340), .B0(n4015), .B1(n6660), .Y(
        n6801) );
  OAI22XL U1720 ( .A0(n7011), .A1(n4008), .B0(n4193), .B1(n4360), .Y(n6660) );
  AOI22X2 U1721 ( .A0(mem_rdata[101]), .A1(n1340), .B0(n4015), .B1(n6661), .Y(
        n6802) );
  OAI22XL U1722 ( .A0(n7016), .A1(n4008), .B0(n4193), .B1(n4361), .Y(n6661) );
  AOI22X2 U1723 ( .A0(mem_rdata[102]), .A1(n1340), .B0(n4010), .B1(n6662), .Y(
        n6803) );
  OAI22XL U1724 ( .A0(n7021), .A1(n4008), .B0(n4193), .B1(n4362), .Y(n6662) );
  AOI22X2 U1725 ( .A0(mem_rdata[103]), .A1(n1340), .B0(n4012), .B1(n6663), .Y(
        n6804) );
  OAI22XL U1726 ( .A0(n7026), .A1(n4008), .B0(n4193), .B1(n4363), .Y(n6663) );
  AOI22X2 U1727 ( .A0(mem_rdata[104]), .A1(n1340), .B0(n4018), .B1(n6664), .Y(
        n6805) );
  OAI22XL U1728 ( .A0(n7031), .A1(n4008), .B0(n4192), .B1(n4364), .Y(n6664) );
  AOI22X2 U1729 ( .A0(mem_rdata[118]), .A1(n1339), .B0(n4016), .B1(n6678), .Y(
        n6819) );
  OAI22XL U1730 ( .A0(n6951), .A1(n4008), .B0(n4192), .B1(n4378), .Y(n6678) );
  AOI22X2 U1731 ( .A0(mem_rdata[119]), .A1(n1339), .B0(n4016), .B1(n6679), .Y(
        n6820) );
  OAI22XL U1732 ( .A0(n6956), .A1(n4008), .B0(n4192), .B1(n4379), .Y(n6679) );
  AOI22X2 U1733 ( .A0(mem_rdata[120]), .A1(n1339), .B0(n4016), .B1(n6680), .Y(
        n6821) );
  OAI22XL U1734 ( .A0(n6961), .A1(n6687), .B0(n4192), .B1(n4380), .Y(n6680) );
  AOI22X2 U1735 ( .A0(mem_rdata[121]), .A1(n1339), .B0(n4016), .B1(n6681), .Y(
        n6822) );
  OAI22XL U1736 ( .A0(n6966), .A1(n6687), .B0(n7036), .B1(n4381), .Y(n6681) );
  AOI22X2 U1737 ( .A0(mem_rdata[122]), .A1(n1338), .B0(n4016), .B1(n6682), .Y(
        n6823) );
  OAI22XL U1738 ( .A0(n6971), .A1(n6687), .B0(n7036), .B1(n4382), .Y(n6682) );
  AOI22X2 U1739 ( .A0(mem_rdata[123]), .A1(n1338), .B0(n4016), .B1(n6683), .Y(
        n6824) );
  OAI22XL U1740 ( .A0(n6976), .A1(n6687), .B0(n7036), .B1(n4383), .Y(n6683) );
  AOI22X2 U1741 ( .A0(mem_rdata[124]), .A1(n1338), .B0(n4016), .B1(n6684), .Y(
        n6825) );
  OAI22XL U1742 ( .A0(n6981), .A1(n6687), .B0(n4192), .B1(n4384), .Y(n6684) );
  AOI22X2 U1743 ( .A0(mem_rdata[125]), .A1(n1338), .B0(n4016), .B1(n6685), .Y(
        n6826) );
  OAI22XL U1744 ( .A0(n6986), .A1(n6687), .B0(n4192), .B1(n4385), .Y(n6685) );
  AOI22X2 U1745 ( .A0(mem_rdata[126]), .A1(n1338), .B0(n4017), .B1(n6686), .Y(
        n6827) );
  OAI22XL U1746 ( .A0(n6996), .A1(n6687), .B0(n4192), .B1(n4386), .Y(n6686) );
  AOI22X2 U1747 ( .A0(mem_rdata[127]), .A1(n1338), .B0(n4017), .B1(n6688), .Y(
        n6828) );
  OAI22XL U1748 ( .A0(n7001), .A1(n6687), .B0(n4192), .B1(n4387), .Y(n6688) );
  AOI22X2 U1749 ( .A0(mem_rdata[0]), .A1(n1338), .B0(n4017), .B1(n6689), .Y(
        n6862) );
  OAI22XL U1750 ( .A0(n7038), .A1(n4356), .B0(n6882), .B1(n4009), .Y(n6689) );
  AOI22X2 U1751 ( .A0(mem_rdata[1]), .A1(n1338), .B0(n4017), .B1(n6690), .Y(
        n6863) );
  OAI22XL U1752 ( .A0(n4195), .A1(n4357), .B0(n6937), .B1(n4009), .Y(n6690) );
  AOI22X2 U1753 ( .A0(mem_rdata[2]), .A1(n1338), .B0(n4017), .B1(n6691), .Y(
        n6864) );
  OAI22XL U1754 ( .A0(n4195), .A1(n4358), .B0(n6992), .B1(n4009), .Y(n6691) );
  AOI22X2 U1755 ( .A0(mem_rdata[3]), .A1(n1338), .B0(n4017), .B1(n6692), .Y(
        n6865) );
  OAI22XL U1756 ( .A0(n4195), .A1(n4359), .B0(n7007), .B1(n4009), .Y(n6692) );
  AOI22X2 U1757 ( .A0(mem_rdata[4]), .A1(n1338), .B0(n4017), .B1(n6693), .Y(
        n6866) );
  OAI22XL U1758 ( .A0(n4195), .A1(n4360), .B0(n7012), .B1(n4009), .Y(n6693) );
  AOI22X2 U1759 ( .A0(mem_rdata[5]), .A1(n1337), .B0(n4017), .B1(n6694), .Y(
        n6867) );
  OAI22XL U1760 ( .A0(n4195), .A1(n4361), .B0(n7017), .B1(n4009), .Y(n6694) );
  AOI22X2 U1761 ( .A0(mem_rdata[18]), .A1(n1345), .B0(n4010), .B1(n6575), .Y(
        n6719) );
  OAI22XL U1762 ( .A0(n4195), .A1(n4374), .B0(n6927), .B1(n6706), .Y(n6575) );
  AOI22X2 U1763 ( .A0(mem_rdata[35]), .A1(n1340), .B0(n4011), .B1(n6592), .Y(
        n6736) );
  OAI22XL U1764 ( .A0(n4199), .A1(n4359), .B0(n7009), .B1(n6620), .Y(n6592) );
  AOI22X2 U1765 ( .A0(mem_rdata[36]), .A1(n1337), .B0(n4011), .B1(n6593), .Y(
        n6737) );
  OAI22XL U1766 ( .A0(n4198), .A1(n4360), .B0(n7014), .B1(n6620), .Y(n6593) );
  AOI22X2 U1767 ( .A0(mem_rdata[37]), .A1(n1341), .B0(n4011), .B1(n6594), .Y(
        n6738) );
  OAI22XL U1768 ( .A0(n4199), .A1(n4361), .B0(n7019), .B1(n6620), .Y(n6594) );
  AOI22X2 U1769 ( .A0(mem_rdata[38]), .A1(n1344), .B0(n4011), .B1(n6595), .Y(
        n6739) );
  OAI22XL U1770 ( .A0(n4198), .A1(n4362), .B0(n7024), .B1(n6620), .Y(n6595) );
  AOI22X2 U1771 ( .A0(mem_rdata[39]), .A1(n1344), .B0(n4011), .B1(n6596), .Y(
        n6740) );
  OAI22XL U1772 ( .A0(n4199), .A1(n4363), .B0(n7029), .B1(n6620), .Y(n6596) );
  AOI22X2 U1773 ( .A0(mem_rdata[40]), .A1(n1344), .B0(n4011), .B1(n6597), .Y(
        n6741) );
  OAI22XL U1774 ( .A0(n4199), .A1(n4364), .B0(n7034), .B1(n4006), .Y(n6597) );
  AOI22X2 U1775 ( .A0(mem_rdata[41]), .A1(n1344), .B0(n4011), .B1(n6598), .Y(
        n6742) );
  OAI22XL U1776 ( .A0(n4199), .A1(n4365), .B0(n7042), .B1(n4006), .Y(n6598) );
  AOI22X2 U1777 ( .A0(mem_rdata[42]), .A1(n1344), .B0(n4012), .B1(n6599), .Y(
        n6743) );
  OAI22XL U1778 ( .A0(n4199), .A1(n4366), .B0(n6889), .B1(n4006), .Y(n6599) );
  AOI22X2 U1779 ( .A0(mem_rdata[43]), .A1(n1344), .B0(n4012), .B1(n6600), .Y(
        n6744) );
  OAI22XL U1780 ( .A0(n4199), .A1(n4367), .B0(n6894), .B1(n4006), .Y(n6600) );
  AOI22X2 U1781 ( .A0(mem_rdata[44]), .A1(n1344), .B0(n4012), .B1(n6601), .Y(
        n6745) );
  OAI22XL U1782 ( .A0(n4198), .A1(n4368), .B0(n6899), .B1(n4006), .Y(n6601) );
  AOI22X2 U1783 ( .A0(mem_rdata[45]), .A1(n1344), .B0(n4012), .B1(n6602), .Y(
        n6746) );
  OAI22XL U1784 ( .A0(n4199), .A1(n4369), .B0(n6904), .B1(n4006), .Y(n6602) );
  AOI22X2 U1785 ( .A0(mem_rdata[46]), .A1(n1344), .B0(n4012), .B1(n6603), .Y(
        n6747) );
  OAI22XL U1786 ( .A0(n4198), .A1(n4370), .B0(n6909), .B1(n4006), .Y(n6603) );
  AOI22X2 U1787 ( .A0(mem_rdata[47]), .A1(n1344), .B0(n4012), .B1(n6604), .Y(
        n6748) );
  OAI22XL U1788 ( .A0(n4199), .A1(n4371), .B0(n6914), .B1(n4006), .Y(n6604) );
  AOI22X2 U1789 ( .A0(mem_rdata[48]), .A1(n1344), .B0(n4012), .B1(n6605), .Y(
        n6749) );
  OAI22XL U1790 ( .A0(n4201), .A1(n4372), .B0(n6919), .B1(n4006), .Y(n6605) );
  AOI22X2 U1791 ( .A0(mem_rdata[49]), .A1(n1344), .B0(n4012), .B1(n6606), .Y(
        n6750) );
  OAI22XL U1792 ( .A0(n4199), .A1(n4373), .B0(n6924), .B1(n4006), .Y(n6606) );
  AOI22X2 U1793 ( .A0(mem_rdata[50]), .A1(n1343), .B0(n4012), .B1(n6607), .Y(
        n6751) );
  OAI22XL U1794 ( .A0(n4199), .A1(n4374), .B0(n6929), .B1(n4006), .Y(n6607) );
  AOI22X2 U1795 ( .A0(mem_rdata[51]), .A1(n1343), .B0(n4012), .B1(n6608), .Y(
        n6752) );
  OAI22XL U1796 ( .A0(n4199), .A1(n4375), .B0(n6934), .B1(n4006), .Y(n6608) );
  AOI22X2 U1797 ( .A0(mem_rdata[52]), .A1(n1343), .B0(n4012), .B1(n6609), .Y(
        n6753) );
  OAI22XL U1798 ( .A0(n4199), .A1(n4376), .B0(n6944), .B1(n4006), .Y(n6609) );
  AOI22X2 U1799 ( .A0(mem_rdata[53]), .A1(n1343), .B0(n4012), .B1(n6610), .Y(
        n6754) );
  OAI22XL U1800 ( .A0(n7041), .A1(n4377), .B0(n6949), .B1(n4006), .Y(n6610) );
  AOI22X2 U1801 ( .A0(mem_rdata[54]), .A1(n1343), .B0(n4013), .B1(n6611), .Y(
        n6755) );
  OAI22XL U1802 ( .A0(n7041), .A1(n4378), .B0(n6954), .B1(n4006), .Y(n6611) );
  AOI22X2 U1803 ( .A0(mem_rdata[55]), .A1(n1343), .B0(n4013), .B1(n6612), .Y(
        n6756) );
  OAI22XL U1804 ( .A0(n7041), .A1(n4379), .B0(n6959), .B1(n4006), .Y(n6612) );
  AOI22X2 U1805 ( .A0(mem_rdata[56]), .A1(n1343), .B0(n4013), .B1(n6613), .Y(
        n6757) );
  OAI22XL U1806 ( .A0(n7041), .A1(n4380), .B0(n6964), .B1(n6620), .Y(n6613) );
  AOI22X2 U1807 ( .A0(mem_rdata[57]), .A1(n1343), .B0(n4013), .B1(n6614), .Y(
        n6758) );
  OAI22XL U1808 ( .A0(n7041), .A1(n4381), .B0(n6969), .B1(n6620), .Y(n6614) );
  AOI22X2 U1809 ( .A0(mem_rdata[58]), .A1(n1343), .B0(n4013), .B1(n6615), .Y(
        n6759) );
  OAI22XL U1810 ( .A0(n4198), .A1(n4382), .B0(n6974), .B1(n6620), .Y(n6615) );
  AOI22X2 U1811 ( .A0(mem_rdata[59]), .A1(n1343), .B0(n4013), .B1(n6616), .Y(
        n6760) );
  OAI22XL U1812 ( .A0(n4199), .A1(n4383), .B0(n6979), .B1(n6620), .Y(n6616) );
  AOI22X2 U1813 ( .A0(mem_rdata[60]), .A1(n1343), .B0(n4013), .B1(n6617), .Y(
        n6761) );
  OAI22XL U1814 ( .A0(n4198), .A1(n4384), .B0(n6984), .B1(n6620), .Y(n6617) );
  AOI22X2 U1815 ( .A0(mem_rdata[61]), .A1(n1343), .B0(n4013), .B1(n6618), .Y(
        n6762) );
  OAI22XL U1816 ( .A0(n4199), .A1(n4385), .B0(n6989), .B1(n6620), .Y(n6618) );
  AOI22X2 U1817 ( .A0(mem_rdata[62]), .A1(n1342), .B0(n4013), .B1(n6619), .Y(
        n6763) );
  OAI22XL U1818 ( .A0(n4198), .A1(n4386), .B0(n6999), .B1(n6620), .Y(n6619) );
  AOI22X2 U1819 ( .A0(mem_rdata[63]), .A1(n1342), .B0(n4013), .B1(n6621), .Y(
        n6764) );
  OAI22XL U1820 ( .A0(n4199), .A1(n4387), .B0(n7004), .B1(n6620), .Y(n6621) );
  AOI22X2 U1821 ( .A0(mem_rdata[64]), .A1(n1342), .B0(n4013), .B1(n6623), .Y(
        n6765) );
  OAI22XL U1822 ( .A0(n4203), .A1(n4356), .B0(n6885), .B1(n6654), .Y(n6623) );
  AOI22X2 U1823 ( .A0(mem_rdata[65]), .A1(n1342), .B0(n4013), .B1(n6624), .Y(
        n6766) );
  OAI22XL U1824 ( .A0(n4203), .A1(n4357), .B0(n6940), .B1(n6654), .Y(n6624) );
  AOI22X2 U1825 ( .A0(mem_rdata[66]), .A1(n1342), .B0(n4014), .B1(n6625), .Y(
        n6767) );
  OAI22XL U1826 ( .A0(n4203), .A1(n4358), .B0(n6995), .B1(n6654), .Y(n6625) );
  AOI22X2 U1827 ( .A0(mem_rdata[67]), .A1(n1342), .B0(n4014), .B1(n6626), .Y(
        n6768) );
  OAI22XL U1828 ( .A0(n4203), .A1(n4359), .B0(n7010), .B1(n6654), .Y(n6626) );
  AOI22X2 U1829 ( .A0(mem_rdata[68]), .A1(n1342), .B0(n4014), .B1(n6627), .Y(
        n6769) );
  OAI22XL U1830 ( .A0(n4203), .A1(n4360), .B0(n7015), .B1(n6654), .Y(n6627) );
  AOI22X2 U1831 ( .A0(mem_rdata[69]), .A1(n1342), .B0(n4014), .B1(n6628), .Y(
        n6770) );
  OAI22XL U1832 ( .A0(n4203), .A1(n4361), .B0(n7020), .B1(n4007), .Y(n6628) );
  AOI22X2 U1833 ( .A0(mem_rdata[70]), .A1(n1342), .B0(n4014), .B1(n6629), .Y(
        n6771) );
  OAI22XL U1834 ( .A0(n4202), .A1(n4362), .B0(n7025), .B1(n4007), .Y(n6629) );
  AOI22X2 U1835 ( .A0(mem_rdata[71]), .A1(n1342), .B0(n4014), .B1(n6630), .Y(
        n6772) );
  OAI22XL U1836 ( .A0(n4203), .A1(n4363), .B0(n7030), .B1(n4007), .Y(n6630) );
  AOI22X2 U1837 ( .A0(mem_rdata[72]), .A1(n1342), .B0(n4014), .B1(n6631), .Y(
        n6773) );
  OAI22XL U1838 ( .A0(n4203), .A1(n4364), .B0(n7035), .B1(n4007), .Y(n6631) );
  AOI22X2 U1839 ( .A0(mem_rdata[73]), .A1(n1342), .B0(n4014), .B1(n6632), .Y(
        n6774) );
  OAI22XL U1840 ( .A0(n4202), .A1(n4365), .B0(n7044), .B1(n4007), .Y(n6632) );
  AOI22X2 U1841 ( .A0(mem_rdata[74]), .A1(n1343), .B0(n4014), .B1(n6633), .Y(
        n6775) );
  OAI22XL U1842 ( .A0(n4202), .A1(n4366), .B0(n6890), .B1(n4007), .Y(n6633) );
  AOI22X2 U1843 ( .A0(mem_rdata[75]), .A1(n1342), .B0(n4014), .B1(n6634), .Y(
        n6776) );
  OAI22XL U1844 ( .A0(n4202), .A1(n4367), .B0(n6895), .B1(n4007), .Y(n6634) );
  AOI22X2 U1845 ( .A0(mem_rdata[76]), .A1(n1340), .B0(n4014), .B1(n6635), .Y(
        n6777) );
  OAI22XL U1846 ( .A0(n4202), .A1(n4368), .B0(n6900), .B1(n4007), .Y(n6635) );
  AOI22X2 U1847 ( .A0(mem_rdata[77]), .A1(n1341), .B0(n4014), .B1(n6636), .Y(
        n6778) );
  OAI22XL U1848 ( .A0(n4203), .A1(n4369), .B0(n6905), .B1(n4007), .Y(n6636) );
  AOI22X2 U1849 ( .A0(mem_rdata[78]), .A1(n1343), .B0(n4011), .B1(n6637), .Y(
        n6779) );
  OAI22XL U1850 ( .A0(n4202), .A1(n4370), .B0(n6910), .B1(n4007), .Y(n6637) );
  AOI22X2 U1851 ( .A0(mem_rdata[79]), .A1(n1342), .B0(n4014), .B1(n6638), .Y(
        n6780) );
  OAI22XL U1852 ( .A0(n4203), .A1(n4371), .B0(n6915), .B1(n4007), .Y(n6638) );
  AOI22X2 U1853 ( .A0(mem_rdata[80]), .A1(n1345), .B0(n4011), .B1(n6639), .Y(
        n6781) );
  OAI22XL U1854 ( .A0(n4202), .A1(n4372), .B0(n6920), .B1(n4007), .Y(n6639) );
  AOI22X2 U1855 ( .A0(mem_rdata[81]), .A1(n1338), .B0(n4017), .B1(n6640), .Y(
        n6782) );
  OAI22XL U1856 ( .A0(n4203), .A1(n4373), .B0(n6925), .B1(n4007), .Y(n6640) );
  AOI22X2 U1857 ( .A0(mem_rdata[82]), .A1(n1338), .B0(n4016), .B1(n6641), .Y(
        n6783) );
  OAI22XL U1858 ( .A0(n4202), .A1(n4374), .B0(n6930), .B1(n4007), .Y(n6641) );
  AOI22X2 U1859 ( .A0(mem_rdata[83]), .A1(n4351), .B0(n4014), .B1(n6642), .Y(
        n6784) );
  OAI22XL U1860 ( .A0(n4203), .A1(n4375), .B0(n6935), .B1(n4007), .Y(n6642) );
  AOI22X2 U1861 ( .A0(mem_rdata[84]), .A1(n4351), .B0(n4017), .B1(n6643), .Y(
        n6785) );
  OAI22XL U1862 ( .A0(n4205), .A1(n4376), .B0(n6945), .B1(n4007), .Y(n6643) );
  AOI22X2 U1863 ( .A0(mem_rdata[85]), .A1(n4351), .B0(n4016), .B1(n6644), .Y(
        n6786) );
  OAI22XL U1864 ( .A0(n4202), .A1(n4377), .B0(n6950), .B1(n4007), .Y(n6644) );
  AOI22X2 U1865 ( .A0(mem_rdata[86]), .A1(n1341), .B0(n4017), .B1(n6645), .Y(
        n6787) );
  OAI22XL U1866 ( .A0(n4202), .A1(n4378), .B0(n6955), .B1(n4007), .Y(n6645) );
  AOI22X2 U1867 ( .A0(mem_rdata[87]), .A1(n1341), .B0(n4016), .B1(n6646), .Y(
        n6788) );
  OAI22XL U1868 ( .A0(n4202), .A1(n4379), .B0(n6960), .B1(n4007), .Y(n6646) );
  AOI22X2 U1869 ( .A0(mem_rdata[88]), .A1(n1341), .B0(n4011), .B1(n6647), .Y(
        n6789) );
  OAI22XL U1870 ( .A0(n4202), .A1(n4380), .B0(n6965), .B1(n6654), .Y(n6647) );
  AOI22X2 U1871 ( .A0(mem_rdata[105]), .A1(n1340), .B0(n4018), .B1(n6665), .Y(
        n6806) );
  OAI22XL U1872 ( .A0(n7037), .A1(n6687), .B0(n4192), .B1(n4365), .Y(n6665) );
  AOI22X2 U1873 ( .A0(mem_rdata[106]), .A1(n1340), .B0(n4018), .B1(n6666), .Y(
        n6807) );
  OAI22XL U1874 ( .A0(n6886), .A1(n6687), .B0(n4192), .B1(n4366), .Y(n6666) );
  AOI22X2 U1875 ( .A0(mem_rdata[107]), .A1(n1340), .B0(n4018), .B1(n6667), .Y(
        n6808) );
  OAI22XL U1876 ( .A0(n6891), .A1(n6687), .B0(n4192), .B1(n4367), .Y(n6667) );
  AOI22X2 U1877 ( .A0(mem_rdata[108]), .A1(n1340), .B0(n4018), .B1(n6668), .Y(
        n6809) );
  OAI22XL U1878 ( .A0(n6896), .A1(n4008), .B0(n4192), .B1(n4368), .Y(n6668) );
  AOI22X2 U1879 ( .A0(mem_rdata[109]), .A1(n1340), .B0(n4013), .B1(n6669), .Y(
        n6810) );
  OAI22XL U1880 ( .A0(n6901), .A1(n4008), .B0(n4192), .B1(n4369), .Y(n6669) );
  AOI22X2 U1881 ( .A0(mem_rdata[110]), .A1(n1339), .B0(n4010), .B1(n6670), .Y(
        n6811) );
  OAI22XL U1882 ( .A0(n6906), .A1(n4008), .B0(n4192), .B1(n4370), .Y(n6670) );
  AOI22X2 U1883 ( .A0(mem_rdata[111]), .A1(n1339), .B0(n4013), .B1(n6671), .Y(
        n6812) );
  OAI22XL U1884 ( .A0(n6911), .A1(n4008), .B0(n4192), .B1(n4371), .Y(n6671) );
  AOI22X2 U1885 ( .A0(mem_rdata[112]), .A1(n1339), .B0(n4012), .B1(n6672), .Y(
        n6813) );
  OAI22XL U1886 ( .A0(n6916), .A1(n4008), .B0(n4192), .B1(n4372), .Y(n6672) );
  AOI22X2 U1887 ( .A0(mem_rdata[113]), .A1(n1339), .B0(n4018), .B1(n6673), .Y(
        n6814) );
  OAI22XL U1888 ( .A0(n6921), .A1(n4008), .B0(n4192), .B1(n4373), .Y(n6673) );
  AOI22X2 U1889 ( .A0(mem_rdata[114]), .A1(n1339), .B0(n4016), .B1(n6674), .Y(
        n6815) );
  OAI22XL U1890 ( .A0(n6926), .A1(n4008), .B0(n4192), .B1(n4374), .Y(n6674) );
  AOI22X2 U1891 ( .A0(mem_rdata[115]), .A1(n1339), .B0(n4016), .B1(n6675), .Y(
        n6816) );
  OAI22XL U1892 ( .A0(n6931), .A1(n4008), .B0(n4192), .B1(n4375), .Y(n6675) );
  AOI22X2 U1893 ( .A0(mem_rdata[116]), .A1(n1339), .B0(n4016), .B1(n6676), .Y(
        n6817) );
  OAI22XL U1894 ( .A0(n6941), .A1(n4008), .B0(n4194), .B1(n4376), .Y(n6676) );
  AOI22X2 U1895 ( .A0(mem_rdata[117]), .A1(n1339), .B0(n4016), .B1(n6677), .Y(
        n6818) );
  OAI22XL U1896 ( .A0(n6946), .A1(n4008), .B0(n4192), .B1(n4377), .Y(n6677) );
  AOI22X2 U1897 ( .A0(mem_rdata[6]), .A1(n1337), .B0(n4017), .B1(n6695), .Y(
        n6868) );
  OAI22XL U1898 ( .A0(n4195), .A1(n4362), .B0(n7022), .B1(n4009), .Y(n6695) );
  AOI22X2 U1899 ( .A0(mem_rdata[7]), .A1(n1337), .B0(n4017), .B1(n6696), .Y(
        n6869) );
  OAI22XL U1900 ( .A0(n4195), .A1(n4363), .B0(n7027), .B1(n4009), .Y(n6696) );
  AOI22X2 U1901 ( .A0(mem_rdata[8]), .A1(n1337), .B0(n4017), .B1(n6697), .Y(
        n6870) );
  OAI22XL U1902 ( .A0(n4195), .A1(n4364), .B0(n7032), .B1(n4009), .Y(n6697) );
  AOI22X2 U1903 ( .A0(mem_rdata[9]), .A1(n1337), .B0(n4017), .B1(n6698), .Y(
        n6871) );
  OAI22XL U1904 ( .A0(n7038), .A1(n4365), .B0(n7039), .B1(n4009), .Y(n6698) );
  AOI22X2 U1905 ( .A0(mem_rdata[10]), .A1(n1337), .B0(n4018), .B1(n6699), .Y(
        n6872) );
  OAI22XL U1906 ( .A0(n4195), .A1(n4366), .B0(n6887), .B1(n6706), .Y(n6699) );
  AOI22X2 U1907 ( .A0(mem_rdata[11]), .A1(n1337), .B0(n4018), .B1(n6700), .Y(
        n6873) );
  OAI22XL U1908 ( .A0(n4195), .A1(n4367), .B0(n6892), .B1(n6706), .Y(n6700) );
  AOI22X2 U1909 ( .A0(mem_rdata[12]), .A1(n1337), .B0(n4018), .B1(n6701), .Y(
        n6874) );
  OAI22XL U1910 ( .A0(n4195), .A1(n4368), .B0(n6897), .B1(n6706), .Y(n6701) );
  AOI22X2 U1911 ( .A0(mem_rdata[13]), .A1(n1337), .B0(n4018), .B1(n6702), .Y(
        n6875) );
  OAI22XL U1912 ( .A0(n7038), .A1(n4369), .B0(n6902), .B1(n6706), .Y(n6702) );
  AOI22X2 U1913 ( .A0(mem_rdata[14]), .A1(n1337), .B0(n4018), .B1(n6703), .Y(
        n6876) );
  OAI22XL U1914 ( .A0(n4195), .A1(n4370), .B0(n6907), .B1(n6706), .Y(n6703) );
  AOI22X2 U1915 ( .A0(mem_rdata[15]), .A1(n1337), .B0(n4018), .B1(n6704), .Y(
        n6877) );
  OAI22XL U1916 ( .A0(n4195), .A1(n4371), .B0(n6912), .B1(n6706), .Y(n6704) );
  AOI22X2 U1917 ( .A0(mem_rdata[16]), .A1(n1337), .B0(n4018), .B1(n6705), .Y(
        n6878) );
  OAI22XL U1918 ( .A0(n4195), .A1(n4372), .B0(n6917), .B1(n6706), .Y(n6705) );
  AOI22X2 U1919 ( .A0(mem_rdata[17]), .A1(n1337), .B0(n4018), .B1(n6707), .Y(
        n6879) );
  OAI22XL U1920 ( .A0(n4195), .A1(n4373), .B0(n6922), .B1(n6706), .Y(n6707) );
  NOR2X1 U1921 ( .A(\state_r[0] ), .B(n8289), .Y(n6832) );
  NAND2X2 U1922 ( .A(\state_r[0] ), .B(n8272), .Y(n7045) );
  OAI22XL U1923 ( .A0(n4137), .A1(n8063), .B0(n4148), .B1(n8191), .Y(n6070) );
  OAI22XL U1924 ( .A0(n4117), .A1(n7807), .B0(n4128), .B1(n7935), .Y(n6069) );
  OAI22XL U1925 ( .A0(n1696), .A1(n7551), .B0(n1355), .B1(n7679), .Y(n6072) );
  OAI22XL U1926 ( .A0(n4137), .A1(n8064), .B0(n4148), .B1(n8192), .Y(n6074) );
  OAI22XL U1927 ( .A0(n4117), .A1(n7808), .B0(n4128), .B1(n7936), .Y(n6073) );
  OAI22XL U1928 ( .A0(n1693), .A1(n7552), .B0(n1356), .B1(n7680), .Y(n6076) );
  OAI22XL U1929 ( .A0(n4137), .A1(n8065), .B0(n4148), .B1(n8193), .Y(n6082) );
  OAI22XL U1930 ( .A0(n4117), .A1(n7809), .B0(n4128), .B1(n7937), .Y(n6081) );
  OAI22XL U1931 ( .A0(n1696), .A1(n7553), .B0(n1357), .B1(n7681), .Y(n6084) );
  OAI22XL U1932 ( .A0(n4137), .A1(n8066), .B0(n4148), .B1(n8194), .Y(n6086) );
  OAI22XL U1933 ( .A0(n4117), .A1(n7810), .B0(n4128), .B1(n7938), .Y(n6085) );
  OAI22XL U1934 ( .A0(n1693), .A1(n7554), .B0(n1354), .B1(n7682), .Y(n6088) );
  OAI22XL U1935 ( .A0(n4137), .A1(n8067), .B0(n4148), .B1(n8195), .Y(n6090) );
  OAI22XL U1936 ( .A0(n4117), .A1(n7811), .B0(n4128), .B1(n7939), .Y(n6089) );
  OAI22XL U1937 ( .A0(n1696), .A1(n7555), .B0(n1356), .B1(n7683), .Y(n6092) );
  OAI22XL U1938 ( .A0(n4137), .A1(n8068), .B0(n4148), .B1(n8196), .Y(n6094) );
  OAI22XL U1939 ( .A0(n4117), .A1(n7812), .B0(n4128), .B1(n7940), .Y(n6093) );
  OAI22XL U1940 ( .A0(n1697), .A1(n7556), .B0(n1357), .B1(n7684), .Y(n6096) );
  OAI22XL U1941 ( .A0(n4137), .A1(n8069), .B0(n4148), .B1(n8197), .Y(n6098) );
  OAI22XL U1942 ( .A0(n4117), .A1(n7813), .B0(n4128), .B1(n7941), .Y(n6097) );
  OAI22XL U1943 ( .A0(n1695), .A1(n7557), .B0(n1355), .B1(n7685), .Y(n6100) );
  OAI22XL U1944 ( .A0(n4137), .A1(n8070), .B0(n4148), .B1(n8198), .Y(n6102) );
  OAI22XL U1945 ( .A0(n4117), .A1(n7814), .B0(n4128), .B1(n7942), .Y(n6101) );
  OAI22XL U1946 ( .A0(n1695), .A1(n7558), .B0(n1354), .B1(n7686), .Y(n6104) );
  OAI22XL U1947 ( .A0(n4137), .A1(n8071), .B0(n4148), .B1(n8199), .Y(n6106) );
  OAI22XL U1948 ( .A0(n4117), .A1(n7815), .B0(n4128), .B1(n7943), .Y(n6105) );
  OAI22XL U1949 ( .A0(n1693), .A1(n7559), .B0(n1354), .B1(n7687), .Y(n6108) );
  OAI22XL U1950 ( .A0(n4137), .A1(n8072), .B0(n4148), .B1(n8200), .Y(n6110) );
  OAI22XL U1951 ( .A0(n4117), .A1(n7816), .B0(n4128), .B1(n7944), .Y(n6109) );
  OAI22XL U1952 ( .A0(n1695), .A1(n7560), .B0(n1356), .B1(n7688), .Y(n6112) );
  OAI22XL U1953 ( .A0(n4136), .A1(n8076), .B0(n4147), .B1(n8204), .Y(n6130) );
  OAI22XL U1954 ( .A0(n4116), .A1(n7820), .B0(n4127), .B1(n7948), .Y(n6129) );
  OAI22XL U1955 ( .A0(n1701), .A1(n7564), .B0(n1358), .B1(n7692), .Y(n6132) );
  OAI22XL U1956 ( .A0(n4136), .A1(n8077), .B0(n4147), .B1(n8205), .Y(n6134) );
  OAI22XL U1957 ( .A0(n4116), .A1(n7821), .B0(n4127), .B1(n7949), .Y(n6133) );
  OAI22XL U1958 ( .A0(n1701), .A1(n7565), .B0(n1358), .B1(n7693), .Y(n6136) );
  OAI22XL U1959 ( .A0(n4136), .A1(n8078), .B0(n4147), .B1(n8206), .Y(n6138) );
  OAI22XL U1960 ( .A0(n4116), .A1(n7822), .B0(n4127), .B1(n7950), .Y(n6137) );
  OAI22XL U1961 ( .A0(n1701), .A1(n7566), .B0(n1358), .B1(n7694), .Y(n6140) );
  OAI22XL U1962 ( .A0(n4136), .A1(n8073), .B0(n4147), .B1(n8201), .Y(n6114) );
  OAI22XL U1963 ( .A0(n4116), .A1(n7817), .B0(n4127), .B1(n7945), .Y(n6113) );
  OAI22XL U1964 ( .A0(n1701), .A1(n7561), .B0(n1358), .B1(n7689), .Y(n6116) );
  OAI22XL U1965 ( .A0(n4141), .A1(n8095), .B0(n4146), .B1(n8223), .Y(n6214) );
  OAI22XL U1966 ( .A0(n4121), .A1(n7839), .B0(n4126), .B1(n7967), .Y(n6213) );
  OAI22XL U1967 ( .A0(n1695), .A1(n7583), .B0(n1357), .B1(n7711), .Y(n6216) );
  OAI22XL U1968 ( .A0(n4141), .A1(n8096), .B0(n4146), .B1(n8224), .Y(n6218) );
  OAI22XL U1969 ( .A0(n4116), .A1(n7840), .B0(n4126), .B1(n7968), .Y(n6217) );
  OAI22XL U1970 ( .A0(n1693), .A1(n7584), .B0(n1357), .B1(n7712), .Y(n6220) );
  OAI22XL U1971 ( .A0(n4136), .A1(n8097), .B0(n4146), .B1(n8225), .Y(n6222) );
  OAI22XL U1972 ( .A0(n4121), .A1(n7841), .B0(n4126), .B1(n7969), .Y(n6221) );
  OAI22XL U1973 ( .A0(n2628), .A1(n7585), .B0(n1355), .B1(n7713), .Y(n6224) );
  OAI22XL U1974 ( .A0(n4138), .A1(n8098), .B0(n4146), .B1(n8226), .Y(n6226) );
  OAI22XL U1975 ( .A0(n4118), .A1(n7842), .B0(n4126), .B1(n7970), .Y(n6225) );
  OAI22XL U1976 ( .A0(n1693), .A1(n7586), .B0(n1357), .B1(n7714), .Y(n6228) );
  OAI22XL U1977 ( .A0(n4138), .A1(n8099), .B0(n4146), .B1(n8227), .Y(n6230) );
  OAI22XL U1978 ( .A0(n4118), .A1(n7843), .B0(n4126), .B1(n7971), .Y(n6229) );
  OAI22XL U1979 ( .A0(n1695), .A1(n7587), .B0(n1357), .B1(n7715), .Y(n6232) );
  OAI22XL U1980 ( .A0(n4138), .A1(n8100), .B0(n4146), .B1(n8228), .Y(n6234) );
  OAI22XL U1981 ( .A0(n4118), .A1(n7844), .B0(n4126), .B1(n7972), .Y(n6233) );
  OAI22XL U1982 ( .A0(n1693), .A1(n7588), .B0(n1357), .B1(n7716), .Y(n6236) );
  OAI22XL U1983 ( .A0(n4136), .A1(n8101), .B0(n4146), .B1(n8229), .Y(n6238) );
  OAI22XL U1984 ( .A0(n4116), .A1(n7845), .B0(n4126), .B1(n7973), .Y(n6237) );
  OAI22XL U1985 ( .A0(n1695), .A1(n7589), .B0(n1357), .B1(n7717), .Y(n6240) );
  OAI22XL U1986 ( .A0(n4141), .A1(n8102), .B0(n4146), .B1(n8230), .Y(n6242) );
  OAI22XL U1987 ( .A0(n4116), .A1(n7846), .B0(n4126), .B1(n7974), .Y(n6241) );
  OAI22XL U1988 ( .A0(n2628), .A1(n7590), .B0(n1358), .B1(n7718), .Y(n6244) );
  OAI22XL U1989 ( .A0(n4136), .A1(n8103), .B0(n4146), .B1(n8231), .Y(n6246) );
  OAI22XL U1990 ( .A0(n4116), .A1(n7847), .B0(n4126), .B1(n7975), .Y(n6245) );
  OAI22XL U1991 ( .A0(n1693), .A1(n7591), .B0(n1355), .B1(n7719), .Y(n6248) );
  OAI22XL U1992 ( .A0(n4135), .A1(n8104), .B0(n4145), .B1(n8232), .Y(n6250) );
  OAI22XL U1993 ( .A0(n4115), .A1(n7848), .B0(n4125), .B1(n7976), .Y(n6249) );
  OAI22XL U1994 ( .A0(n1697), .A1(n7592), .B0(n1580), .B1(n7720), .Y(n6252) );
  OAI22XL U1995 ( .A0(n4135), .A1(n8108), .B0(n4145), .B1(n8236), .Y(n6270) );
  OAI22XL U1996 ( .A0(n4115), .A1(n7852), .B0(n4125), .B1(n7980), .Y(n6269) );
  OAI22XL U1997 ( .A0(n1697), .A1(n7596), .B0(n1354), .B1(n7724), .Y(n6272) );
  OAI22XL U1998 ( .A0(n4135), .A1(n8109), .B0(n4145), .B1(n8237), .Y(n6274) );
  OAI22XL U1999 ( .A0(n4115), .A1(n7853), .B0(n4125), .B1(n7981), .Y(n6273) );
  OAI22XL U2000 ( .A0(n1697), .A1(n7597), .B0(n1355), .B1(n7725), .Y(n6276) );
  OAI22XL U2001 ( .A0(n4135), .A1(n8110), .B0(n4145), .B1(n8238), .Y(n6278) );
  OAI22XL U2002 ( .A0(n4115), .A1(n7854), .B0(n4125), .B1(n7982), .Y(n6277) );
  OAI22XL U2003 ( .A0(n1697), .A1(n7598), .B0(n1354), .B1(n7726), .Y(n6280) );
  OAI22XL U2004 ( .A0(n4135), .A1(n8105), .B0(n4145), .B1(n8233), .Y(n6258) );
  OAI22XL U2005 ( .A0(n4115), .A1(n7849), .B0(n4125), .B1(n7977), .Y(n6257) );
  OAI22XL U2006 ( .A0(n1697), .A1(n7593), .B0(n1356), .B1(n7721), .Y(n6260) );
  OAI22XL U2007 ( .A0(n4140), .A1(n8127), .B0(n4144), .B1(n8255), .Y(n5846) );
  OAI22XL U2008 ( .A0(n4120), .A1(n7871), .B0(n6846), .B1(n7999), .Y(n5845) );
  OAI22XL U2009 ( .A0(n1696), .A1(n7615), .B0(n1357), .B1(n7743), .Y(n5848) );
  OAI22XL U2010 ( .A0(n4140), .A1(n8128), .B0(n6849), .B1(n8256), .Y(n5850) );
  OAI22XL U2011 ( .A0(n4120), .A1(n7872), .B0(n6846), .B1(n8000), .Y(n5849) );
  OAI22XL U2012 ( .A0(n1697), .A1(n7616), .B0(n1355), .B1(n7744), .Y(n5852) );
  OAI22XL U2013 ( .A0(n4140), .A1(n8129), .B0(n6849), .B1(n8257), .Y(n5854) );
  OAI22XL U2014 ( .A0(n4120), .A1(n7873), .B0(n6846), .B1(n8001), .Y(n5853) );
  OAI22XL U2015 ( .A0(n1695), .A1(n7617), .B0(n1356), .B1(n7745), .Y(n5856) );
  OAI22XL U2016 ( .A0(n4140), .A1(n8130), .B0(n4144), .B1(n8258), .Y(n5858) );
  OAI22XL U2017 ( .A0(n4120), .A1(n7874), .B0(n4125), .B1(n8002), .Y(n5857) );
  OAI22XL U2018 ( .A0(n1704), .A1(n7618), .B0(n1354), .B1(n7746), .Y(n5860) );
  OAI22XL U2019 ( .A0(n4140), .A1(n8131), .B0(n4144), .B1(n8259), .Y(n5862) );
  OAI22XL U2020 ( .A0(n4120), .A1(n7875), .B0(n4130), .B1(n8003), .Y(n5861) );
  OAI22XL U2021 ( .A0(n1696), .A1(n7619), .B0(n1357), .B1(n7747), .Y(n5864) );
  OAI22XL U2022 ( .A0(n4140), .A1(n8132), .B0(n4144), .B1(n8260), .Y(n5866) );
  OAI22XL U2023 ( .A0(n4120), .A1(n7876), .B0(n4124), .B1(n8004), .Y(n5865) );
  OAI22XL U2024 ( .A0(n1693), .A1(n7620), .B0(n1355), .B1(n7748), .Y(n5868) );
  OAI22XL U2025 ( .A0(n4140), .A1(n8133), .B0(n6849), .B1(n8261), .Y(n5870) );
  OAI22XL U2026 ( .A0(n4120), .A1(n7877), .B0(n4124), .B1(n8005), .Y(n5869) );
  OAI22XL U2027 ( .A0(n1703), .A1(n7621), .B0(n1356), .B1(n7749), .Y(n5872) );
  OAI22XL U2028 ( .A0(n4140), .A1(n8134), .B0(n6849), .B1(n8262), .Y(n5874) );
  OAI22XL U2029 ( .A0(n4120), .A1(n7878), .B0(n4124), .B1(n8006), .Y(n5873) );
  OAI22XL U2030 ( .A0(n1704), .A1(n7622), .B0(n1354), .B1(n7750), .Y(n5876) );
  OAI22XL U2031 ( .A0(n4140), .A1(n8135), .B0(n6849), .B1(n8263), .Y(n5882) );
  OAI22XL U2032 ( .A0(n4120), .A1(n7879), .B0(n6846), .B1(n8007), .Y(n5881) );
  OAI22XL U2033 ( .A0(n1696), .A1(n7623), .B0(n1354), .B1(n7751), .Y(n5884) );
  OAI22XL U2034 ( .A0(n4140), .A1(n8136), .B0(n6849), .B1(n8264), .Y(n5886) );
  OAI22XL U2035 ( .A0(n4120), .A1(n7880), .B0(n6846), .B1(n8008), .Y(n5885) );
  OAI22XL U2036 ( .A0(n1693), .A1(n7624), .B0(n1357), .B1(n7752), .Y(n5888) );
  OAI22XL U2037 ( .A0(n4140), .A1(n8137), .B0(n4144), .B1(n8265), .Y(n5890) );
  OAI22XL U2038 ( .A0(n4120), .A1(n7881), .B0(n6846), .B1(n8009), .Y(n5889) );
  OAI22XL U2039 ( .A0(n1695), .A1(n7625), .B0(n1355), .B1(n7753), .Y(n5892) );
  OAI22XL U2040 ( .A0(n4140), .A1(n8140), .B0(n4150), .B1(n8268), .Y(n5902) );
  OAI22XL U2041 ( .A0(n4120), .A1(n7884), .B0(n4125), .B1(n8012), .Y(n5901) );
  OAI22XL U2042 ( .A0(n1696), .A1(n7628), .B0(n1357), .B1(n7756), .Y(n5904) );
  OAI22XL U2043 ( .A0(n4140), .A1(n8141), .B0(n4150), .B1(n8269), .Y(n5906) );
  OAI22XL U2044 ( .A0(n4120), .A1(n7885), .B0(n4131), .B1(n8013), .Y(n5905) );
  OAI22XL U2045 ( .A0(n1693), .A1(n7629), .B0(n1528), .B1(n7757), .Y(n5908) );
  OAI22XL U2046 ( .A0(n4140), .A1(n8142), .B0(n4151), .B1(n8270), .Y(n5910) );
  OAI22XL U2047 ( .A0(n4120), .A1(n7886), .B0(n4130), .B1(n8014), .Y(n5909) );
  OAI22XL U2048 ( .A0(n1701), .A1(n7630), .B0(n1355), .B1(n7758), .Y(n5912) );
  OAI22XL U2049 ( .A0(n4139), .A1(n8033), .B0(n4150), .B1(n8161), .Y(n5938) );
  OAI22XL U2050 ( .A0(n4119), .A1(n7777), .B0(n4130), .B1(n7905), .Y(n5937) );
  OAI22XL U2051 ( .A0(n1704), .A1(n7521), .B0(n1528), .B1(n7649), .Y(n5940) );
  OAI22XL U2052 ( .A0(n4139), .A1(n8034), .B0(n4150), .B1(n8162), .Y(n5942) );
  OAI22XL U2053 ( .A0(n4119), .A1(n7778), .B0(n4130), .B1(n7906), .Y(n5941) );
  OAI22XL U2054 ( .A0(n1704), .A1(n7522), .B0(n1528), .B1(n7650), .Y(n5944) );
  OAI22XL U2055 ( .A0(n4139), .A1(n8035), .B0(n4150), .B1(n8163), .Y(n5950) );
  OAI22XL U2056 ( .A0(n4119), .A1(n7779), .B0(n4130), .B1(n7907), .Y(n5949) );
  OAI22XL U2057 ( .A0(n1704), .A1(n7523), .B0(n1528), .B1(n7651), .Y(n5952) );
  OAI22XL U2058 ( .A0(n4139), .A1(n8036), .B0(n4150), .B1(n8164), .Y(n5954) );
  OAI22XL U2059 ( .A0(n4119), .A1(n7780), .B0(n4130), .B1(n7908), .Y(n5953) );
  OAI22XL U2060 ( .A0(n1704), .A1(n7524), .B0(n1528), .B1(n7652), .Y(n5956) );
  OAI22XL U2061 ( .A0(n4139), .A1(n8037), .B0(n4150), .B1(n8165), .Y(n5958) );
  OAI22XL U2062 ( .A0(n4119), .A1(n7781), .B0(n4130), .B1(n7909), .Y(n5957) );
  OAI22XL U2063 ( .A0(n1704), .A1(n7525), .B0(n1528), .B1(n7653), .Y(n5960) );
  OAI22XL U2064 ( .A0(n4139), .A1(n8038), .B0(n4150), .B1(n8166), .Y(n5962) );
  OAI22XL U2065 ( .A0(n4119), .A1(n7782), .B0(n4130), .B1(n7910), .Y(n5961) );
  OAI22XL U2066 ( .A0(n1704), .A1(n7526), .B0(n1528), .B1(n7654), .Y(n5964) );
  OAI22XL U2067 ( .A0(n4139), .A1(n8039), .B0(n4150), .B1(n8167), .Y(n5966) );
  OAI22XL U2068 ( .A0(n4119), .A1(n7783), .B0(n4130), .B1(n7911), .Y(n5965) );
  OAI22XL U2069 ( .A0(n1704), .A1(n7527), .B0(n1528), .B1(n7655), .Y(n5968) );
  OAI22XL U2070 ( .A0(n4139), .A1(n8040), .B0(n4150), .B1(n8168), .Y(n5970) );
  OAI22XL U2071 ( .A0(n4119), .A1(n7784), .B0(n4130), .B1(n7912), .Y(n5969) );
  OAI22XL U2072 ( .A0(n1704), .A1(n7528), .B0(n1528), .B1(n7656), .Y(n5972) );
  OAI22XL U2073 ( .A0(n4139), .A1(n8041), .B0(n4150), .B1(n8169), .Y(n5974) );
  OAI22XL U2074 ( .A0(n4119), .A1(n7785), .B0(n4130), .B1(n7913), .Y(n5973) );
  OAI22XL U2075 ( .A0(n1704), .A1(n7529), .B0(n1528), .B1(n7657), .Y(n5976) );
  OAI22XL U2076 ( .A0(n4138), .A1(n8044), .B0(n4149), .B1(n8172), .Y(n5986) );
  OAI22XL U2077 ( .A0(n4118), .A1(n7788), .B0(n4129), .B1(n7916), .Y(n5985) );
  OAI22XL U2078 ( .A0(n1703), .A1(n7532), .B0(n1359), .B1(n7660), .Y(n5988) );
  OAI22XL U2079 ( .A0(n4138), .A1(n8045), .B0(n4149), .B1(n8173), .Y(n5994) );
  OAI22XL U2080 ( .A0(n4118), .A1(n7789), .B0(n4129), .B1(n7917), .Y(n5993) );
  OAI22XL U2081 ( .A0(n1703), .A1(n7533), .B0(n1359), .B1(n7661), .Y(n5996) );
  OAI22XL U2082 ( .A0(n4138), .A1(n8046), .B0(n4149), .B1(n8174), .Y(n5998) );
  OAI22XL U2083 ( .A0(n4118), .A1(n7790), .B0(n4129), .B1(n7918), .Y(n5997) );
  OAI22XL U2084 ( .A0(n1703), .A1(n7534), .B0(n1359), .B1(n7662), .Y(n6000) );
  OAI22XL U2085 ( .A0(n4139), .A1(n8031), .B0(n4150), .B1(n8159), .Y(n5930) );
  OAI22XL U2086 ( .A0(n4119), .A1(n7775), .B0(n4130), .B1(n7903), .Y(n5929) );
  OAI22XL U2087 ( .A0(n1704), .A1(n7519), .B0(n1528), .B1(n7647), .Y(n5932) );
  OAI22XL U2088 ( .A0(n4139), .A1(n8032), .B0(n4150), .B1(n8160), .Y(n5934) );
  OAI22XL U2089 ( .A0(n4119), .A1(n7776), .B0(n4130), .B1(n7904), .Y(n5933) );
  OAI22XL U2090 ( .A0(n1704), .A1(n7520), .B0(n1528), .B1(n7648), .Y(n5936) );
  OAI32X1 U2091 ( .A0(n6837), .A1(n4352), .A2(n6840), .B0(n6842), .B1(n8272), 
        .Y(n4423) );
  OAI22XL U2092 ( .A0(n4040), .A1(n7522), .B0(n6720), .B1(n4036), .Y(n4915) );
  OAI22XL U2093 ( .A0(n4054), .A1(n7650), .B0(n6720), .B1(n4051), .Y(n5043) );
  OAI22XL U2094 ( .A0(n4083), .A1(n7906), .B0(n6720), .B1(n4080), .Y(n5299) );
  OAI22XL U2095 ( .A0(n4094), .A1(n8034), .B0(n6720), .B1(n4087), .Y(n5427) );
  OAI22XL U2096 ( .A0(n4108), .A1(n8162), .B0(n6720), .B1(n4101), .Y(n5555) );
  OAI22XL U2097 ( .A0(n4187), .A1(n7266), .B0(n6720), .B1(n4178), .Y(n4659) );
  OAI22XL U2098 ( .A0(n4040), .A1(n7523), .B0(n6721), .B1(n4036), .Y(n4916) );
  OAI22XL U2099 ( .A0(n4054), .A1(n7651), .B0(n6721), .B1(n4051), .Y(n5044) );
  OAI22XL U2100 ( .A0(n4083), .A1(n7907), .B0(n6721), .B1(n4080), .Y(n5300) );
  OAI22XL U2101 ( .A0(n4094), .A1(n8035), .B0(n6721), .B1(n4087), .Y(n5428) );
  OAI22XL U2102 ( .A0(n4108), .A1(n8163), .B0(n6721), .B1(n4101), .Y(n5556) );
  OAI22XL U2103 ( .A0(n4186), .A1(n7267), .B0(n6721), .B1(n4178), .Y(n4660) );
  OAI22XL U2104 ( .A0(n4040), .A1(n7524), .B0(n6722), .B1(n4032), .Y(n4917) );
  OAI22XL U2105 ( .A0(n4056), .A1(n7652), .B0(n6722), .B1(n4046), .Y(n5045) );
  OAI22XL U2106 ( .A0(n4083), .A1(n7908), .B0(n6722), .B1(n4080), .Y(n5301) );
  OAI22XL U2107 ( .A0(n4094), .A1(n8036), .B0(n6722), .B1(n4087), .Y(n5429) );
  OAI22XL U2108 ( .A0(n4108), .A1(n8164), .B0(n6722), .B1(n4101), .Y(n5557) );
  OAI22XL U2109 ( .A0(n4185), .A1(n7268), .B0(n6722), .B1(n4178), .Y(n4661) );
  OAI22XL U2110 ( .A0(n4040), .A1(n7525), .B0(n6723), .B1(n4037), .Y(n4918) );
  OAI22XL U2111 ( .A0(n4055), .A1(n7653), .B0(n6723), .B1(n4050), .Y(n5046) );
  OAI22XL U2112 ( .A0(n4083), .A1(n7909), .B0(n6723), .B1(n4080), .Y(n5302) );
  OAI22XL U2113 ( .A0(n4094), .A1(n8037), .B0(n6723), .B1(n4087), .Y(n5430) );
  OAI22XL U2114 ( .A0(n4108), .A1(n8165), .B0(n6723), .B1(n4101), .Y(n5558) );
  OAI22XL U2115 ( .A0(n4189), .A1(n7269), .B0(n6723), .B1(n4178), .Y(n4662) );
  OAI22XL U2116 ( .A0(n4040), .A1(n7526), .B0(n6724), .B1(n4035), .Y(n4919) );
  OAI22XL U2117 ( .A0(n4056), .A1(n7654), .B0(n6724), .B1(n4049), .Y(n5047) );
  OAI22XL U2118 ( .A0(n4083), .A1(n7910), .B0(n6724), .B1(n4080), .Y(n5303) );
  OAI22XL U2119 ( .A0(n4094), .A1(n8038), .B0(n6724), .B1(n4087), .Y(n5431) );
  OAI22XL U2120 ( .A0(n4108), .A1(n8166), .B0(n6724), .B1(n4101), .Y(n5559) );
  OAI22XL U2121 ( .A0(n4187), .A1(n7270), .B0(n6724), .B1(n4178), .Y(n4663) );
  OAI22XL U2122 ( .A0(n4041), .A1(n7527), .B0(n6725), .B1(n4032), .Y(n4920) );
  OAI22XL U2123 ( .A0(n4058), .A1(n7655), .B0(n6725), .B1(n4046), .Y(n5048) );
  OAI22XL U2124 ( .A0(n4083), .A1(n7911), .B0(n6725), .B1(n4080), .Y(n5304) );
  OAI22XL U2125 ( .A0(n4095), .A1(n8039), .B0(n6725), .B1(n4088), .Y(n5432) );
  OAI22XL U2126 ( .A0(n4109), .A1(n8167), .B0(n6725), .B1(n4102), .Y(n5560) );
  OAI22XL U2127 ( .A0(n4186), .A1(n7271), .B0(n6725), .B1(n4178), .Y(n4664) );
  OAI22XL U2128 ( .A0(n4041), .A1(n7528), .B0(n6726), .B1(n4032), .Y(n4921) );
  OAI22XL U2129 ( .A0(n4058), .A1(n7656), .B0(n6726), .B1(n4046), .Y(n5049) );
  OAI22XL U2130 ( .A0(n4083), .A1(n7912), .B0(n6726), .B1(n4080), .Y(n5305) );
  OAI22XL U2131 ( .A0(n4095), .A1(n8040), .B0(n6726), .B1(n4088), .Y(n5433) );
  OAI22XL U2132 ( .A0(n4109), .A1(n8168), .B0(n6726), .B1(n4102), .Y(n5561) );
  OAI22XL U2133 ( .A0(n4185), .A1(n7272), .B0(n6726), .B1(n4178), .Y(n4665) );
  OAI22XL U2134 ( .A0(n4041), .A1(n7529), .B0(n6727), .B1(n4032), .Y(n4922) );
  OAI22XL U2135 ( .A0(n4058), .A1(n7657), .B0(n6727), .B1(n4046), .Y(n5050) );
  OAI22XL U2136 ( .A0(n4083), .A1(n7913), .B0(n6727), .B1(n4080), .Y(n5306) );
  OAI22XL U2137 ( .A0(n4095), .A1(n8041), .B0(n6727), .B1(n4088), .Y(n5434) );
  OAI22XL U2138 ( .A0(n4109), .A1(n8169), .B0(n6727), .B1(n4102), .Y(n5562) );
  OAI22XL U2139 ( .A0(n4190), .A1(n7273), .B0(n6727), .B1(n4178), .Y(n4666) );
  OAI22XL U2140 ( .A0(n4041), .A1(n7530), .B0(n6728), .B1(n4032), .Y(n4923) );
  OAI22XL U2141 ( .A0(n4058), .A1(n7658), .B0(n6728), .B1(n4046), .Y(n5051) );
  OAI22XL U2142 ( .A0(n4083), .A1(n7914), .B0(n6728), .B1(n4080), .Y(n5307) );
  OAI22XL U2143 ( .A0(n4095), .A1(n8042), .B0(n6728), .B1(n4088), .Y(n5435) );
  OAI22XL U2144 ( .A0(n4109), .A1(n8170), .B0(n6728), .B1(n4102), .Y(n5563) );
  OAI22XL U2145 ( .A0(n4189), .A1(n7274), .B0(n6728), .B1(n4178), .Y(n4667) );
  OAI22XL U2146 ( .A0(n4041), .A1(n7531), .B0(n6729), .B1(n4032), .Y(n4924) );
  OAI22XL U2147 ( .A0(n4058), .A1(n7659), .B0(n6729), .B1(n4046), .Y(n5052) );
  OAI22XL U2148 ( .A0(n4083), .A1(n7915), .B0(n6729), .B1(n4080), .Y(n5308) );
  OAI22XL U2149 ( .A0(n4095), .A1(n8043), .B0(n6729), .B1(n4088), .Y(n5436) );
  OAI22XL U2150 ( .A0(n4109), .A1(n8171), .B0(n6729), .B1(n4102), .Y(n5564) );
  OAI22XL U2151 ( .A0(n4187), .A1(n7275), .B0(n6729), .B1(n4178), .Y(n4668) );
  OAI22XL U2152 ( .A0(n4041), .A1(n7532), .B0(n6730), .B1(n4032), .Y(n4925) );
  OAI22XL U2153 ( .A0(n4058), .A1(n7660), .B0(n6730), .B1(n4046), .Y(n5053) );
  OAI22XL U2154 ( .A0(n4083), .A1(n7916), .B0(n6730), .B1(n4080), .Y(n5309) );
  OAI22XL U2155 ( .A0(n4095), .A1(n8044), .B0(n6730), .B1(n4088), .Y(n5437) );
  OAI22XL U2156 ( .A0(n4109), .A1(n8172), .B0(n6730), .B1(n4102), .Y(n5565) );
  OAI22XL U2157 ( .A0(n4186), .A1(n7276), .B0(n6730), .B1(n4178), .Y(n4669) );
  OAI22XL U2158 ( .A0(n4041), .A1(n7533), .B0(n6731), .B1(n4032), .Y(n4926) );
  OAI22XL U2159 ( .A0(n4058), .A1(n7661), .B0(n6731), .B1(n4046), .Y(n5054) );
  OAI22XL U2160 ( .A0(n4084), .A1(n7917), .B0(n6731), .B1(n4080), .Y(n5310) );
  OAI22XL U2161 ( .A0(n4095), .A1(n8045), .B0(n6731), .B1(n4088), .Y(n5438) );
  OAI22XL U2162 ( .A0(n4109), .A1(n8173), .B0(n6731), .B1(n4102), .Y(n5566) );
  OAI22XL U2163 ( .A0(n4190), .A1(n7277), .B0(n6731), .B1(n4183), .Y(n4670) );
  OAI22XL U2164 ( .A0(n4041), .A1(n7534), .B0(n6732), .B1(n4032), .Y(n4927) );
  OAI22XL U2165 ( .A0(n4055), .A1(n7662), .B0(n6732), .B1(n4046), .Y(n5055) );
  OAI22XL U2166 ( .A0(n4084), .A1(n7918), .B0(n6732), .B1(n4080), .Y(n5311) );
  OAI22XL U2167 ( .A0(n4095), .A1(n8046), .B0(n6732), .B1(n4088), .Y(n5439) );
  OAI22XL U2168 ( .A0(n4109), .A1(n8174), .B0(n6732), .B1(n4102), .Y(n5567) );
  OAI22XL U2169 ( .A0(n4185), .A1(n7278), .B0(n6732), .B1(n4183), .Y(n4671) );
  OAI22XL U2170 ( .A0(n4041), .A1(n7535), .B0(n6733), .B1(n4032), .Y(n4928) );
  OAI22XL U2171 ( .A0(n4054), .A1(n7663), .B0(n6733), .B1(n4046), .Y(n5056) );
  OAI22XL U2172 ( .A0(n4084), .A1(n7919), .B0(n6733), .B1(n4079), .Y(n5312) );
  OAI22XL U2173 ( .A0(n4095), .A1(n8047), .B0(n6733), .B1(n4088), .Y(n5440) );
  OAI22XL U2174 ( .A0(n4109), .A1(n8175), .B0(n6733), .B1(n4102), .Y(n5568) );
  OAI22XL U2175 ( .A0(n4190), .A1(n7279), .B0(n6733), .B1(n4183), .Y(n4672) );
  OAI22XL U2176 ( .A0(n4041), .A1(n7536), .B0(n6734), .B1(n4032), .Y(n4929) );
  OAI22XL U2177 ( .A0(n4056), .A1(n7664), .B0(n6734), .B1(n4046), .Y(n5057) );
  OAI22XL U2178 ( .A0(n4084), .A1(n7920), .B0(n6734), .B1(n4079), .Y(n5313) );
  OAI22XL U2179 ( .A0(n4095), .A1(n8048), .B0(n6734), .B1(n4088), .Y(n5441) );
  OAI22XL U2180 ( .A0(n4109), .A1(n8176), .B0(n6734), .B1(n4102), .Y(n5569) );
  OAI22XL U2181 ( .A0(n4185), .A1(n7280), .B0(n6734), .B1(n4183), .Y(n4673) );
  OAI22XL U2182 ( .A0(n4041), .A1(n7537), .B0(n6735), .B1(n4032), .Y(n4930) );
  OAI22XL U2183 ( .A0(n4056), .A1(n7665), .B0(n6735), .B1(n4046), .Y(n5058) );
  OAI22XL U2184 ( .A0(n4084), .A1(n7921), .B0(n6735), .B1(n4079), .Y(n5314) );
  OAI22XL U2185 ( .A0(n4095), .A1(n8049), .B0(n6735), .B1(n4088), .Y(n5442) );
  OAI22XL U2186 ( .A0(n4109), .A1(n8177), .B0(n6735), .B1(n4102), .Y(n5570) );
  OAI22XL U2187 ( .A0(n4188), .A1(n7281), .B0(n6735), .B1(n4183), .Y(n4674) );
  OAI22XL U2188 ( .A0(n4043), .A1(n7592), .B0(n6790), .B1(n4037), .Y(n4985) );
  OAI22XL U2189 ( .A0(n4056), .A1(n7720), .B0(n6790), .B1(n4050), .Y(n5113) );
  OAI22XL U2190 ( .A0(n4065), .A1(n7848), .B0(n6790), .B1(n4070), .Y(n5241) );
  OAI22XL U2191 ( .A0(n4095), .A1(n8104), .B0(n6790), .B1(n4092), .Y(n5497) );
  OAI22XL U2192 ( .A0(n4109), .A1(n8232), .B0(n6790), .B1(n4106), .Y(n5625) );
  OAI22XL U2193 ( .A0(n4186), .A1(n7336), .B0(n6790), .B1(n4181), .Y(n4729) );
  OAI22XL U2194 ( .A0(n4039), .A1(n7593), .B0(n6791), .B1(n4037), .Y(n4986) );
  OAI22XL U2195 ( .A0(n4056), .A1(n7721), .B0(n6791), .B1(n4050), .Y(n5114) );
  OAI22XL U2196 ( .A0(n4065), .A1(n7849), .B0(n6791), .B1(n4070), .Y(n5242) );
  OAI22XL U2197 ( .A0(n4099), .A1(n8105), .B0(n6791), .B1(n4086), .Y(n5498) );
  OAI22XL U2198 ( .A0(n4113), .A1(n8233), .B0(n6791), .B1(n4100), .Y(n5626) );
  OAI22XL U2199 ( .A0(n4188), .A1(n7337), .B0(n6791), .B1(n4182), .Y(n4730) );
  OAI22XL U2200 ( .A0(n4041), .A1(n7594), .B0(n6792), .B1(n4037), .Y(n4987) );
  OAI22XL U2201 ( .A0(n4056), .A1(n7722), .B0(n6792), .B1(n4050), .Y(n5115) );
  OAI22XL U2202 ( .A0(n4065), .A1(n7850), .B0(n6792), .B1(n4070), .Y(n5243) );
  OAI22XL U2203 ( .A0(n4098), .A1(n8106), .B0(n6792), .B1(n4092), .Y(n5499) );
  OAI22XL U2204 ( .A0(n4112), .A1(n8234), .B0(n6792), .B1(n4106), .Y(n5627) );
  OAI22XL U2205 ( .A0(n4188), .A1(n7338), .B0(n6792), .B1(n4182), .Y(n4731) );
  OAI22XL U2206 ( .A0(n4044), .A1(n7595), .B0(n6793), .B1(n4037), .Y(n4988) );
  OAI22XL U2207 ( .A0(n4056), .A1(n7723), .B0(n6793), .B1(n4050), .Y(n5116) );
  OAI22XL U2208 ( .A0(n4065), .A1(n7851), .B0(n6793), .B1(n4070), .Y(n5244) );
  OAI22XL U2209 ( .A0(n4096), .A1(n8107), .B0(n6793), .B1(n4086), .Y(n5500) );
  OAI22XL U2210 ( .A0(n4110), .A1(n8235), .B0(n6793), .B1(n4100), .Y(n5628) );
  OAI22XL U2211 ( .A0(n4188), .A1(n7339), .B0(n6793), .B1(n4182), .Y(n4732) );
  OAI22XL U2212 ( .A0(n4042), .A1(n7596), .B0(n6794), .B1(n4037), .Y(n4989) );
  OAI22XL U2213 ( .A0(n4056), .A1(n7724), .B0(n6794), .B1(n4050), .Y(n5117) );
  OAI22XL U2214 ( .A0(n4065), .A1(n7852), .B0(n6794), .B1(n4070), .Y(n5245) );
  OAI22XL U2215 ( .A0(n4097), .A1(n8108), .B0(n6794), .B1(n4088), .Y(n5501) );
  OAI22XL U2216 ( .A0(n4111), .A1(n8236), .B0(n6794), .B1(n4102), .Y(n5629) );
  OAI22XL U2217 ( .A0(n4188), .A1(n7340), .B0(n6794), .B1(n4182), .Y(n4733) );
  OAI22XL U2218 ( .A0(n4043), .A1(n7597), .B0(n6795), .B1(n4037), .Y(n4990) );
  OAI22XL U2219 ( .A0(n4056), .A1(n7725), .B0(n6795), .B1(n4050), .Y(n5118) );
  OAI22XL U2220 ( .A0(n4065), .A1(n7853), .B0(n6795), .B1(n4069), .Y(n5246) );
  OAI22XL U2221 ( .A0(n4093), .A1(n8109), .B0(n6795), .B1(n4091), .Y(n5502) );
  OAI22XL U2222 ( .A0(n4107), .A1(n8237), .B0(n6795), .B1(n4105), .Y(n5630) );
  OAI22XL U2223 ( .A0(n4188), .A1(n7341), .B0(n6795), .B1(n4178), .Y(n4734) );
  OAI22XL U2224 ( .A0(n4045), .A1(n7598), .B0(n6796), .B1(n4037), .Y(n4991) );
  OAI22XL U2225 ( .A0(n4056), .A1(n7726), .B0(n6796), .B1(n4050), .Y(n5119) );
  OAI22XL U2226 ( .A0(n4065), .A1(n7854), .B0(n6796), .B1(n4071), .Y(n5247) );
  OAI22XL U2227 ( .A0(n4094), .A1(n8110), .B0(n6796), .B1(n4089), .Y(n5503) );
  OAI22XL U2228 ( .A0(n4108), .A1(n8238), .B0(n6796), .B1(n4103), .Y(n5631) );
  OAI22XL U2229 ( .A0(n4188), .A1(n7342), .B0(n6796), .B1(n4181), .Y(n4735) );
  OAI22XL U2230 ( .A0(n4045), .A1(n7503), .B0(n6862), .B1(n4034), .Y(n4896) );
  OAI22XL U2231 ( .A0(n4058), .A1(n7631), .B0(n6862), .B1(n4048), .Y(n5024) );
  OAI22XL U2232 ( .A0(n4065), .A1(n7759), .B0(n6862), .B1(n4068), .Y(n5152) );
  OAI22XL U2233 ( .A0(n4093), .A1(n8015), .B0(n6862), .B1(n4086), .Y(n5408) );
  OAI22XL U2234 ( .A0(n4107), .A1(n8143), .B0(n6862), .B1(n4100), .Y(n5536) );
  OAI22XL U2235 ( .A0(n4188), .A1(n7247), .B0(n6862), .B1(n4184), .Y(n4640) );
  OAI22XL U2236 ( .A0(n4045), .A1(n7504), .B0(n6863), .B1(n4036), .Y(n4897) );
  OAI22XL U2237 ( .A0(n4058), .A1(n7632), .B0(n6863), .B1(n4047), .Y(n5025) );
  OAI22XL U2238 ( .A0(n4064), .A1(n7760), .B0(n6863), .B1(n4073), .Y(n5153) );
  OAI22XL U2239 ( .A0(n4093), .A1(n8016), .B0(n6863), .B1(n4086), .Y(n5409) );
  OAI22XL U2240 ( .A0(n4107), .A1(n8144), .B0(n6863), .B1(n4100), .Y(n5537) );
  OAI22XL U2241 ( .A0(n4189), .A1(n7248), .B0(n6863), .B1(n4184), .Y(n4641) );
  OAI22XL U2242 ( .A0(n4045), .A1(n7505), .B0(n6864), .B1(n4032), .Y(n4898) );
  OAI22XL U2243 ( .A0(n4058), .A1(n7633), .B0(n6864), .B1(n4046), .Y(n5026) );
  OAI22XL U2244 ( .A0(n4060), .A1(n7761), .B0(n6864), .B1(n4073), .Y(n5154) );
  OAI22XL U2245 ( .A0(n4093), .A1(n8017), .B0(n6864), .B1(n4086), .Y(n5410) );
  OAI22XL U2246 ( .A0(n4107), .A1(n8145), .B0(n6864), .B1(n4100), .Y(n5538) );
  OAI22XL U2247 ( .A0(n4187), .A1(n7249), .B0(n6864), .B1(n4184), .Y(n4642) );
  OAI22XL U2248 ( .A0(n4045), .A1(n7506), .B0(n6865), .B1(n4037), .Y(n4899) );
  OAI22XL U2249 ( .A0(n4058), .A1(n7634), .B0(n6865), .B1(n4049), .Y(n5027) );
  OAI22XL U2250 ( .A0(n4060), .A1(n7762), .B0(n6865), .B1(n4073), .Y(n5155) );
  OAI22XL U2251 ( .A0(n4093), .A1(n8018), .B0(n6865), .B1(n4086), .Y(n5411) );
  OAI22XL U2252 ( .A0(n4107), .A1(n8146), .B0(n6865), .B1(n4100), .Y(n5539) );
  OAI22XL U2253 ( .A0(n4186), .A1(n7250), .B0(n6865), .B1(n4184), .Y(n4643) );
  OAI22XL U2254 ( .A0(n4039), .A1(n7507), .B0(n6866), .B1(n4035), .Y(n4900) );
  OAI22XL U2255 ( .A0(n4053), .A1(n7635), .B0(n6866), .B1(n4051), .Y(n5028) );
  OAI22XL U2256 ( .A0(n4065), .A1(n7763), .B0(n6866), .B1(n4073), .Y(n5156) );
  OAI22XL U2257 ( .A0(n4093), .A1(n8019), .B0(n6866), .B1(n4086), .Y(n5412) );
  OAI22XL U2258 ( .A0(n4107), .A1(n8147), .B0(n6866), .B1(n4100), .Y(n5540) );
  OAI22XL U2259 ( .A0(n4187), .A1(n7251), .B0(n6866), .B1(n4184), .Y(n4644) );
  OAI22XL U2260 ( .A0(n4045), .A1(n7508), .B0(n6867), .B1(n4038), .Y(n4901) );
  OAI22XL U2261 ( .A0(n4058), .A1(n7636), .B0(n6867), .B1(n4050), .Y(n5029) );
  OAI22XL U2262 ( .A0(n4061), .A1(n7764), .B0(n6867), .B1(n4073), .Y(n5157) );
  OAI22XL U2263 ( .A0(n4093), .A1(n8020), .B0(n6867), .B1(n4086), .Y(n5413) );
  OAI22XL U2264 ( .A0(n4107), .A1(n8148), .B0(n6867), .B1(n4100), .Y(n5541) );
  OAI22XL U2265 ( .A0(n4190), .A1(n7252), .B0(n6867), .B1(n4184), .Y(n4645) );
  OAI22XL U2266 ( .A0(n4042), .A1(n7599), .B0(n6797), .B1(n4037), .Y(n4992) );
  OAI22XL U2267 ( .A0(n4057), .A1(n7727), .B0(n6797), .B1(n4051), .Y(n5120) );
  OAI22XL U2268 ( .A0(n4065), .A1(n7855), .B0(n6797), .B1(n4069), .Y(n5248) );
  OAI22XL U2269 ( .A0(n4093), .A1(n8111), .B0(n6797), .B1(n4092), .Y(n5504) );
  OAI22XL U2270 ( .A0(n4107), .A1(n8239), .B0(n6797), .B1(n4106), .Y(n5632) );
  OAI22XL U2271 ( .A0(n4188), .A1(n7343), .B0(n6797), .B1(n4181), .Y(n4736) );
  OAI22XL U2272 ( .A0(n4044), .A1(n7600), .B0(n6798), .B1(n4035), .Y(n4993) );
  OAI22XL U2273 ( .A0(n4057), .A1(n7728), .B0(n6798), .B1(n4051), .Y(n5121) );
  OAI22XL U2274 ( .A0(n4065), .A1(n7856), .B0(n6798), .B1(n4069), .Y(n5249) );
  OAI22XL U2275 ( .A0(n4094), .A1(n8112), .B0(n6798), .B1(n4086), .Y(n5505) );
  OAI22XL U2276 ( .A0(n4108), .A1(n8240), .B0(n6798), .B1(n4100), .Y(n5633) );
  OAI22XL U2277 ( .A0(n4188), .A1(n7344), .B0(n6798), .B1(n4179), .Y(n4737) );
  OAI22XL U2278 ( .A0(n4043), .A1(n7601), .B0(n6799), .B1(n4036), .Y(n4994) );
  OAI22XL U2279 ( .A0(n4057), .A1(n7729), .B0(n6799), .B1(n4051), .Y(n5122) );
  OAI22XL U2280 ( .A0(n4065), .A1(n7857), .B0(n6799), .B1(n4069), .Y(n5250) );
  OAI22XL U2281 ( .A0(n4096), .A1(n8113), .B0(n6799), .B1(n4092), .Y(n5506) );
  OAI22XL U2282 ( .A0(n4110), .A1(n8241), .B0(n6799), .B1(n4106), .Y(n5634) );
  OAI22XL U2283 ( .A0(n4188), .A1(n7345), .B0(n6799), .B1(n4180), .Y(n4738) );
  OAI22XL U2284 ( .A0(n4045), .A1(n7602), .B0(n6800), .B1(n4032), .Y(n4995) );
  OAI22XL U2285 ( .A0(n4057), .A1(n7730), .B0(n6800), .B1(n4051), .Y(n5123) );
  OAI22XL U2286 ( .A0(n4065), .A1(n7858), .B0(n6800), .B1(n4069), .Y(n5251) );
  OAI22XL U2287 ( .A0(n4093), .A1(n8114), .B0(n6800), .B1(n4086), .Y(n5507) );
  OAI22XL U2288 ( .A0(n4107), .A1(n8242), .B0(n6800), .B1(n4100), .Y(n5635) );
  OAI22XL U2289 ( .A0(n4188), .A1(n7346), .B0(n6800), .B1(n4181), .Y(n4739) );
  OAI22XL U2290 ( .A0(n4041), .A1(n7603), .B0(n6801), .B1(n4037), .Y(n4996) );
  OAI22XL U2291 ( .A0(n4057), .A1(n7731), .B0(n6801), .B1(n4051), .Y(n5124) );
  OAI22XL U2292 ( .A0(n4065), .A1(n7859), .B0(n6801), .B1(n4069), .Y(n5252) );
  OAI22XL U2293 ( .A0(n4094), .A1(n8115), .B0(n6801), .B1(n4092), .Y(n5508) );
  OAI22XL U2294 ( .A0(n4108), .A1(n8243), .B0(n6801), .B1(n4106), .Y(n5636) );
  OAI22XL U2295 ( .A0(n4188), .A1(n7347), .B0(n6801), .B1(n1), .Y(n4740) );
  OAI22XL U2296 ( .A0(n4042), .A1(n7604), .B0(n6802), .B1(n4035), .Y(n4997) );
  OAI22XL U2297 ( .A0(n4057), .A1(n7732), .B0(n6802), .B1(n4051), .Y(n5125) );
  OAI22XL U2298 ( .A0(n4061), .A1(n7860), .B0(n6802), .B1(n4069), .Y(n5253) );
  OAI22XL U2299 ( .A0(n4099), .A1(n8116), .B0(n6802), .B1(n4086), .Y(n5509) );
  OAI22XL U2300 ( .A0(n4113), .A1(n8244), .B0(n6802), .B1(n4100), .Y(n5637) );
  OAI22XL U2301 ( .A0(n4188), .A1(n7348), .B0(n6802), .B1(n4180), .Y(n4741) );
  OAI22XL U2302 ( .A0(n4041), .A1(n7605), .B0(n6803), .B1(n4038), .Y(n4998) );
  OAI22XL U2303 ( .A0(n4057), .A1(n7733), .B0(n6803), .B1(n4051), .Y(n5126) );
  OAI22XL U2304 ( .A0(n4062), .A1(n7861), .B0(n6803), .B1(n4069), .Y(n5254) );
  OAI22XL U2305 ( .A0(n4099), .A1(n8117), .B0(n6803), .B1(n4092), .Y(n5510) );
  OAI22XL U2306 ( .A0(n4113), .A1(n8245), .B0(n6803), .B1(n4106), .Y(n5638) );
  OAI22XL U2307 ( .A0(n4189), .A1(n7349), .B0(n6803), .B1(n4182), .Y(n4742) );
  OAI22XL U2308 ( .A0(n4044), .A1(n7606), .B0(n6804), .B1(n4038), .Y(n4999) );
  OAI22XL U2309 ( .A0(n4057), .A1(n7734), .B0(n6804), .B1(n4051), .Y(n5127) );
  OAI22XL U2310 ( .A0(n4063), .A1(n7862), .B0(n6804), .B1(n4069), .Y(n5255) );
  OAI22XL U2311 ( .A0(n4099), .A1(n8118), .B0(n6804), .B1(n4086), .Y(n5511) );
  OAI22XL U2312 ( .A0(n4113), .A1(n8246), .B0(n6804), .B1(n4100), .Y(n5639) );
  OAI22XL U2313 ( .A0(n4189), .A1(n7350), .B0(n6804), .B1(n4182), .Y(n4743) );
  OAI22XL U2314 ( .A0(n4042), .A1(n7607), .B0(n6805), .B1(n4038), .Y(n5000) );
  OAI22XL U2315 ( .A0(n4057), .A1(n7735), .B0(n6805), .B1(n4051), .Y(n5128) );
  OAI22XL U2316 ( .A0(n4064), .A1(n7863), .B0(n6805), .B1(n4069), .Y(n5256) );
  OAI22XL U2317 ( .A0(n4099), .A1(n8119), .B0(n6805), .B1(n4092), .Y(n5512) );
  OAI22XL U2318 ( .A0(n4113), .A1(n8247), .B0(n6805), .B1(n4106), .Y(n5640) );
  OAI22XL U2319 ( .A0(n4189), .A1(n7351), .B0(n6805), .B1(n4182), .Y(n4744) );
  OAI22XL U2320 ( .A0(n4040), .A1(n7621), .B0(n6819), .B1(n4033), .Y(n5014) );
  OAI22XL U2321 ( .A0(n4059), .A1(n7749), .B0(n6819), .B1(n4048), .Y(n5142) );
  OAI22XL U2322 ( .A0(n4085), .A1(n8005), .B0(n6819), .B1(n4075), .Y(n5398) );
  OAI22XL U2323 ( .A0(n4095), .A1(n8133), .B0(n6819), .B1(n4092), .Y(n5526) );
  OAI22XL U2324 ( .A0(n4109), .A1(n8261), .B0(n6819), .B1(n4106), .Y(n5654) );
  OAI22XL U2325 ( .A0(n4190), .A1(n7365), .B0(n6819), .B1(n4183), .Y(n4758) );
  OAI22XL U2326 ( .A0(n4040), .A1(n7622), .B0(n6820), .B1(n4033), .Y(n5015) );
  OAI22XL U2327 ( .A0(n4056), .A1(n7750), .B0(n6820), .B1(n4047), .Y(n5143) );
  OAI22XL U2328 ( .A0(n4082), .A1(n8006), .B0(n6820), .B1(n4075), .Y(n5399) );
  OAI22XL U2329 ( .A0(n4098), .A1(n8134), .B0(n6820), .B1(n4092), .Y(n5527) );
  OAI22XL U2330 ( .A0(n4112), .A1(n8262), .B0(n6820), .B1(n4106), .Y(n5655) );
  OAI22XL U2331 ( .A0(n4190), .A1(n7366), .B0(n6820), .B1(n4183), .Y(n4759) );
  OAI22XL U2332 ( .A0(n4045), .A1(n7623), .B0(n6821), .B1(n4033), .Y(n5016) );
  OAI22XL U2333 ( .A0(n4058), .A1(n7751), .B0(n6821), .B1(n4046), .Y(n5144) );
  OAI22XL U2334 ( .A0(n4083), .A1(n8007), .B0(n6821), .B1(n4074), .Y(n5400) );
  OAI22XL U2335 ( .A0(n4098), .A1(n8135), .B0(n6821), .B1(n4086), .Y(n5528) );
  OAI22XL U2336 ( .A0(n4112), .A1(n8263), .B0(n6821), .B1(n4100), .Y(n5656) );
  OAI22XL U2337 ( .A0(n4190), .A1(n7367), .B0(n6821), .B1(n4183), .Y(n4760) );
  OAI22XL U2338 ( .A0(n4045), .A1(n7624), .B0(n6822), .B1(n4034), .Y(n5017) );
  OAI22XL U2339 ( .A0(n4058), .A1(n7752), .B0(n6822), .B1(n4048), .Y(n5145) );
  OAI22XL U2340 ( .A0(n4082), .A1(n8008), .B0(n6822), .B1(n4075), .Y(n5401) );
  OAI22XL U2341 ( .A0(n4097), .A1(n8136), .B0(n6822), .B1(n4092), .Y(n5529) );
  OAI22XL U2342 ( .A0(n4111), .A1(n8264), .B0(n6822), .B1(n4106), .Y(n5657) );
  OAI22XL U2343 ( .A0(n4190), .A1(n7368), .B0(n6822), .B1(n4183), .Y(n4761) );
  OAI22XL U2344 ( .A0(n4045), .A1(n7625), .B0(n6823), .B1(n5), .Y(n5018) );
  OAI22XL U2345 ( .A0(n4058), .A1(n7753), .B0(n6823), .B1(n6), .Y(n5146) );
  OAI22XL U2346 ( .A0(n4083), .A1(n8009), .B0(n6823), .B1(n4075), .Y(n5402) );
  OAI22XL U2347 ( .A0(n6716), .A1(n8137), .B0(n6823), .B1(n3), .Y(n5530) );
  OAI22XL U2348 ( .A0(n6829), .A1(n8265), .B0(n6823), .B1(n4), .Y(n5658) );
  OAI22XL U2349 ( .A0(n4190), .A1(n7369), .B0(n6823), .B1(n4183), .Y(n4762) );
  OAI22XL U2350 ( .A0(n4045), .A1(n7626), .B0(n6824), .B1(n5), .Y(n5019) );
  OAI22XL U2351 ( .A0(n4058), .A1(n7754), .B0(n6824), .B1(n6), .Y(n5147) );
  OAI22XL U2352 ( .A0(n4081), .A1(n8010), .B0(n6824), .B1(n4075), .Y(n5403) );
  OAI22XL U2353 ( .A0(n4099), .A1(n8138), .B0(n6824), .B1(n3), .Y(n5531) );
  OAI22XL U2354 ( .A0(n4113), .A1(n8266), .B0(n6824), .B1(n4), .Y(n5659) );
  OAI22XL U2355 ( .A0(n4190), .A1(n7370), .B0(n6824), .B1(n4183), .Y(n4763) );
  OAI22XL U2356 ( .A0(n4045), .A1(n7627), .B0(n6825), .B1(n5), .Y(n5020) );
  OAI22XL U2357 ( .A0(n4058), .A1(n7755), .B0(n6825), .B1(n6), .Y(n5148) );
  OAI22XL U2358 ( .A0(n4082), .A1(n8011), .B0(n6825), .B1(n4074), .Y(n5404) );
  OAI22XL U2359 ( .A0(n6716), .A1(n8139), .B0(n6825), .B1(n3), .Y(n5532) );
  OAI22XL U2360 ( .A0(n6829), .A1(n8267), .B0(n6825), .B1(n4), .Y(n5660) );
  OAI22XL U2361 ( .A0(n4190), .A1(n7371), .B0(n6825), .B1(n4183), .Y(n4764) );
  OAI22XL U2362 ( .A0(n4045), .A1(n7628), .B0(n6826), .B1(n5), .Y(n5021) );
  OAI22XL U2363 ( .A0(n4058), .A1(n7756), .B0(n6826), .B1(n6), .Y(n5149) );
  OAI22XL U2364 ( .A0(n4081), .A1(n8012), .B0(n6826), .B1(n4075), .Y(n5405) );
  OAI22XL U2365 ( .A0(n4099), .A1(n8140), .B0(n6826), .B1(n3), .Y(n5533) );
  OAI22XL U2366 ( .A0(n4113), .A1(n8268), .B0(n6826), .B1(n4), .Y(n5661) );
  OAI22XL U2367 ( .A0(n4190), .A1(n7372), .B0(n6826), .B1(n4183), .Y(n4765) );
  OAI22XL U2368 ( .A0(n4045), .A1(n7629), .B0(n6827), .B1(n4033), .Y(n5022) );
  OAI22XL U2369 ( .A0(n4058), .A1(n7757), .B0(n6827), .B1(n4047), .Y(n5150) );
  OAI22XL U2370 ( .A0(n4084), .A1(n8013), .B0(n6827), .B1(n4074), .Y(n5406) );
  OAI22XL U2371 ( .A0(n6716), .A1(n8141), .B0(n6827), .B1(n4089), .Y(n5534) );
  OAI22XL U2372 ( .A0(n6829), .A1(n8269), .B0(n6827), .B1(n4103), .Y(n5662) );
  OAI22XL U2373 ( .A0(n4189), .A1(n7373), .B0(n6827), .B1(n4184), .Y(n4766) );
  OAI22XL U2374 ( .A0(n4045), .A1(n7630), .B0(n6828), .B1(n4034), .Y(n5023) );
  OAI22XL U2375 ( .A0(n4058), .A1(n7758), .B0(n6828), .B1(n4048), .Y(n5151) );
  OAI22XL U2376 ( .A0(n4081), .A1(n8014), .B0(n6828), .B1(n4077), .Y(n5407) );
  OAI22XL U2377 ( .A0(n4099), .A1(n8142), .B0(n6828), .B1(n4090), .Y(n5535) );
  OAI22XL U2378 ( .A0(n4113), .A1(n8270), .B0(n6828), .B1(n4104), .Y(n5663) );
  OAI22XL U2379 ( .A0(n4190), .A1(n7374), .B0(n6828), .B1(n4184), .Y(n4767) );
  OAI22XL U2380 ( .A0(n4040), .A1(n7521), .B0(n6719), .B1(n4036), .Y(n4914) );
  OAI22XL U2381 ( .A0(n4057), .A1(n7649), .B0(n6719), .B1(n4050), .Y(n5042) );
  OAI22XL U2382 ( .A0(n4062), .A1(n7777), .B0(n6719), .B1(n4071), .Y(n5170) );
  OAI22XL U2383 ( .A0(n4083), .A1(n7905), .B0(n6719), .B1(n4074), .Y(n5298) );
  OAI22XL U2384 ( .A0(n4094), .A1(n8033), .B0(n6719), .B1(n4087), .Y(n5426) );
  OAI22XL U2385 ( .A0(n4108), .A1(n8161), .B0(n6719), .B1(n4101), .Y(n5554) );
  OAI22XL U2386 ( .A0(n4185), .A1(n7265), .B0(n6719), .B1(n4178), .Y(n4658) );
  OAI22XL U2387 ( .A0(n4041), .A1(n7538), .B0(n6736), .B1(n4032), .Y(n4931) );
  OAI22XL U2388 ( .A0(n4057), .A1(n7666), .B0(n6736), .B1(n4046), .Y(n5059) );
  OAI22XL U2389 ( .A0(n4063), .A1(n7794), .B0(n6736), .B1(n4071), .Y(n5187) );
  OAI22XL U2390 ( .A0(n4084), .A1(n7922), .B0(n6736), .B1(n4079), .Y(n5315) );
  OAI22XL U2391 ( .A0(n4095), .A1(n8050), .B0(n6736), .B1(n4088), .Y(n5443) );
  OAI22XL U2392 ( .A0(n4109), .A1(n8178), .B0(n6736), .B1(n4102), .Y(n5571) );
  OAI22XL U2393 ( .A0(n4190), .A1(n7282), .B0(n6736), .B1(n4178), .Y(n4675) );
  OAI22XL U2394 ( .A0(n4042), .A1(n7539), .B0(n6737), .B1(n4033), .Y(n4932) );
  OAI22XL U2395 ( .A0(n4054), .A1(n7667), .B0(n6737), .B1(n4047), .Y(n5060) );
  OAI22XL U2396 ( .A0(n4060), .A1(n7795), .B0(n6737), .B1(n4071), .Y(n5188) );
  OAI22XL U2397 ( .A0(n4084), .A1(n7923), .B0(n6737), .B1(n4079), .Y(n5316) );
  OAI22XL U2398 ( .A0(n4096), .A1(n8051), .B0(n6737), .B1(n4089), .Y(n5444) );
  OAI22XL U2399 ( .A0(n4110), .A1(n8179), .B0(n6737), .B1(n4103), .Y(n5572) );
  OAI22XL U2400 ( .A0(n4185), .A1(n7283), .B0(n6737), .B1(n4179), .Y(n4676) );
  OAI22XL U2401 ( .A0(n4042), .A1(n7540), .B0(n6738), .B1(n4033), .Y(n4933) );
  OAI22XL U2402 ( .A0(n4054), .A1(n7668), .B0(n6738), .B1(n4047), .Y(n5061) );
  OAI22XL U2403 ( .A0(n4060), .A1(n7796), .B0(n6738), .B1(n4071), .Y(n5189) );
  OAI22XL U2404 ( .A0(n4084), .A1(n7924), .B0(n6738), .B1(n4079), .Y(n5317) );
  OAI22XL U2405 ( .A0(n4096), .A1(n8052), .B0(n6738), .B1(n4089), .Y(n5445) );
  OAI22XL U2406 ( .A0(n4110), .A1(n8180), .B0(n6738), .B1(n4103), .Y(n5573) );
  OAI22XL U2407 ( .A0(n4188), .A1(n7284), .B0(n6738), .B1(n4181), .Y(n4677) );
  OAI22XL U2408 ( .A0(n4042), .A1(n7541), .B0(n6739), .B1(n4033), .Y(n4934) );
  OAI22XL U2409 ( .A0(n4054), .A1(n7669), .B0(n6739), .B1(n4047), .Y(n5062) );
  OAI22XL U2410 ( .A0(n4060), .A1(n7797), .B0(n6739), .B1(n4071), .Y(n5190) );
  OAI22XL U2411 ( .A0(n4084), .A1(n7925), .B0(n6739), .B1(n4079), .Y(n5318) );
  OAI22XL U2412 ( .A0(n4096), .A1(n8053), .B0(n6739), .B1(n4089), .Y(n5446) );
  OAI22XL U2413 ( .A0(n4110), .A1(n8181), .B0(n6739), .B1(n4103), .Y(n5574) );
  OAI22XL U2414 ( .A0(n4191), .A1(n7285), .B0(n6739), .B1(n4180), .Y(n4678) );
  OAI22XL U2415 ( .A0(n4042), .A1(n7542), .B0(n6740), .B1(n4033), .Y(n4935) );
  OAI22XL U2416 ( .A0(n4054), .A1(n7670), .B0(n6740), .B1(n4047), .Y(n5063) );
  OAI22XL U2417 ( .A0(n4060), .A1(n7798), .B0(n6740), .B1(n4071), .Y(n5191) );
  OAI22XL U2418 ( .A0(n4084), .A1(n7926), .B0(n6740), .B1(n4079), .Y(n5319) );
  OAI22XL U2419 ( .A0(n4096), .A1(n8054), .B0(n6740), .B1(n4089), .Y(n5447) );
  OAI22XL U2420 ( .A0(n4110), .A1(n8182), .B0(n6740), .B1(n4103), .Y(n5575) );
  OAI22XL U2421 ( .A0(n4188), .A1(n7286), .B0(n6740), .B1(n4182), .Y(n4679) );
  OAI22XL U2422 ( .A0(n4042), .A1(n7543), .B0(n6741), .B1(n4033), .Y(n4936) );
  OAI22XL U2423 ( .A0(n4054), .A1(n7671), .B0(n6741), .B1(n4047), .Y(n5064) );
  OAI22XL U2424 ( .A0(n4061), .A1(n7799), .B0(n6741), .B1(n4073), .Y(n5192) );
  OAI22XL U2425 ( .A0(n4084), .A1(n7927), .B0(n6741), .B1(n4079), .Y(n5320) );
  OAI22XL U2426 ( .A0(n4096), .A1(n8055), .B0(n6741), .B1(n4089), .Y(n5448) );
  OAI22XL U2427 ( .A0(n4110), .A1(n8183), .B0(n6741), .B1(n4103), .Y(n5576) );
  OAI22XL U2428 ( .A0(n4191), .A1(n7287), .B0(n6741), .B1(n4184), .Y(n4680) );
  OAI22XL U2429 ( .A0(n4042), .A1(n7544), .B0(n6742), .B1(n4033), .Y(n4937) );
  OAI22XL U2430 ( .A0(n4054), .A1(n7672), .B0(n6742), .B1(n4047), .Y(n5065) );
  OAI22XL U2431 ( .A0(n4061), .A1(n7800), .B0(n6742), .B1(n4070), .Y(n5193) );
  OAI22XL U2432 ( .A0(n4084), .A1(n7928), .B0(n6742), .B1(n4079), .Y(n5321) );
  OAI22XL U2433 ( .A0(n4096), .A1(n8056), .B0(n6742), .B1(n4089), .Y(n5449) );
  OAI22XL U2434 ( .A0(n4110), .A1(n8184), .B0(n6742), .B1(n4103), .Y(n5577) );
  OAI22XL U2435 ( .A0(n4189), .A1(n7288), .B0(n6742), .B1(n4181), .Y(n4681) );
  OAI22XL U2436 ( .A0(n4042), .A1(n7545), .B0(n6743), .B1(n4033), .Y(n4938) );
  OAI22XL U2437 ( .A0(n4054), .A1(n7673), .B0(n6743), .B1(n4047), .Y(n5066) );
  OAI22XL U2438 ( .A0(n4061), .A1(n7801), .B0(n6743), .B1(n4070), .Y(n5194) );
  OAI22XL U2439 ( .A0(n4085), .A1(n7929), .B0(n6743), .B1(n4079), .Y(n5322) );
  OAI22XL U2440 ( .A0(n4096), .A1(n8057), .B0(n6743), .B1(n4089), .Y(n5450) );
  OAI22XL U2441 ( .A0(n4110), .A1(n8185), .B0(n6743), .B1(n4103), .Y(n5578) );
  OAI22XL U2442 ( .A0(n4185), .A1(n7289), .B0(n6743), .B1(n4179), .Y(n4682) );
  OAI22XL U2443 ( .A0(n4042), .A1(n7546), .B0(n6744), .B1(n4033), .Y(n4939) );
  OAI22XL U2444 ( .A0(n4054), .A1(n7674), .B0(n6744), .B1(n4047), .Y(n5067) );
  OAI22XL U2445 ( .A0(n4061), .A1(n7802), .B0(n6744), .B1(n4072), .Y(n5195) );
  OAI22XL U2446 ( .A0(n4085), .A1(n7930), .B0(n6744), .B1(n4079), .Y(n5323) );
  OAI22XL U2447 ( .A0(n4096), .A1(n8058), .B0(n6744), .B1(n4089), .Y(n5451) );
  OAI22XL U2448 ( .A0(n4110), .A1(n8186), .B0(n6744), .B1(n4103), .Y(n5579) );
  OAI22XL U2449 ( .A0(n4185), .A1(n7290), .B0(n6744), .B1(n4179), .Y(n4683) );
  OAI22XL U2450 ( .A0(n4042), .A1(n7547), .B0(n6745), .B1(n4033), .Y(n4940) );
  OAI22XL U2451 ( .A0(n4054), .A1(n7675), .B0(n6745), .B1(n4047), .Y(n5068) );
  OAI22XL U2452 ( .A0(n4061), .A1(n7803), .B0(n6745), .B1(n4072), .Y(n5196) );
  OAI22XL U2453 ( .A0(n4085), .A1(n7931), .B0(n6745), .B1(n4079), .Y(n5324) );
  OAI22XL U2454 ( .A0(n4096), .A1(n8059), .B0(n6745), .B1(n4089), .Y(n5452) );
  OAI22XL U2455 ( .A0(n4110), .A1(n8187), .B0(n6745), .B1(n4103), .Y(n5580) );
  OAI22XL U2456 ( .A0(n4185), .A1(n7291), .B0(n6745), .B1(n4179), .Y(n4684) );
  OAI22XL U2457 ( .A0(n4042), .A1(n7548), .B0(n6746), .B1(n4033), .Y(n4941) );
  OAI22XL U2458 ( .A0(n4054), .A1(n7676), .B0(n6746), .B1(n4047), .Y(n5069) );
  OAI22XL U2459 ( .A0(n4061), .A1(n7804), .B0(n6746), .B1(n4072), .Y(n5197) );
  OAI22XL U2460 ( .A0(n4085), .A1(n7932), .B0(n6746), .B1(n4078), .Y(n5325) );
  OAI22XL U2461 ( .A0(n4096), .A1(n8060), .B0(n6746), .B1(n4089), .Y(n5453) );
  OAI22XL U2462 ( .A0(n4110), .A1(n8188), .B0(n6746), .B1(n4103), .Y(n5581) );
  OAI22XL U2463 ( .A0(n4185), .A1(n7292), .B0(n6746), .B1(n4179), .Y(n4685) );
  OAI22XL U2464 ( .A0(n4042), .A1(n7549), .B0(n6747), .B1(n4033), .Y(n4942) );
  OAI22XL U2465 ( .A0(n4054), .A1(n7677), .B0(n6747), .B1(n4047), .Y(n5070) );
  OAI22XL U2466 ( .A0(n4061), .A1(n7805), .B0(n6747), .B1(n4072), .Y(n5198) );
  OAI22XL U2467 ( .A0(n4085), .A1(n7933), .B0(n6747), .B1(n4078), .Y(n5326) );
  OAI22XL U2468 ( .A0(n4096), .A1(n8061), .B0(n6747), .B1(n4089), .Y(n5454) );
  OAI22XL U2469 ( .A0(n4110), .A1(n8189), .B0(n6747), .B1(n4103), .Y(n5582) );
  OAI22XL U2470 ( .A0(n4185), .A1(n7293), .B0(n6747), .B1(n4179), .Y(n4686) );
  OAI22XL U2471 ( .A0(n4042), .A1(n7550), .B0(n6748), .B1(n4033), .Y(n4943) );
  OAI22XL U2472 ( .A0(n4054), .A1(n7678), .B0(n6748), .B1(n4047), .Y(n5071) );
  OAI22XL U2473 ( .A0(n4061), .A1(n7806), .B0(n6748), .B1(n4072), .Y(n5199) );
  OAI22XL U2474 ( .A0(n4085), .A1(n7934), .B0(n6748), .B1(n4078), .Y(n5327) );
  OAI22XL U2475 ( .A0(n4096), .A1(n8062), .B0(n6748), .B1(n4089), .Y(n5455) );
  OAI22XL U2476 ( .A0(n4110), .A1(n8190), .B0(n6748), .B1(n4103), .Y(n5583) );
  OAI22XL U2477 ( .A0(n4185), .A1(n7294), .B0(n6748), .B1(n4179), .Y(n4687) );
  OAI22XL U2478 ( .A0(n4043), .A1(n7551), .B0(n6749), .B1(n4034), .Y(n4944) );
  OAI22XL U2479 ( .A0(n4059), .A1(n7679), .B0(n6749), .B1(n4048), .Y(n5072) );
  OAI22XL U2480 ( .A0(n4061), .A1(n7807), .B0(n6749), .B1(n4072), .Y(n5200) );
  OAI22XL U2481 ( .A0(n4085), .A1(n7935), .B0(n6749), .B1(n4078), .Y(n5328) );
  OAI22XL U2482 ( .A0(n4097), .A1(n8063), .B0(n6749), .B1(n4090), .Y(n5456) );
  OAI22XL U2483 ( .A0(n4111), .A1(n8191), .B0(n6749), .B1(n4104), .Y(n5584) );
  OAI22XL U2484 ( .A0(n4185), .A1(n7295), .B0(n6749), .B1(n4179), .Y(n4688) );
  OAI22XL U2485 ( .A0(n4043), .A1(n7552), .B0(n6750), .B1(n4034), .Y(n4945) );
  OAI22XL U2486 ( .A0(n4059), .A1(n7680), .B0(n6750), .B1(n4048), .Y(n5073) );
  OAI22XL U2487 ( .A0(n4061), .A1(n7808), .B0(n6750), .B1(n4072), .Y(n5201) );
  OAI22XL U2488 ( .A0(n4085), .A1(n7936), .B0(n6750), .B1(n4078), .Y(n5329) );
  OAI22XL U2489 ( .A0(n4097), .A1(n8064), .B0(n6750), .B1(n4090), .Y(n5457) );
  OAI22XL U2490 ( .A0(n4111), .A1(n8192), .B0(n6750), .B1(n4104), .Y(n5585) );
  OAI22XL U2491 ( .A0(n4185), .A1(n7296), .B0(n6750), .B1(n4179), .Y(n4689) );
  OAI22XL U2492 ( .A0(n4043), .A1(n7553), .B0(n6751), .B1(n4034), .Y(n4946) );
  OAI22XL U2493 ( .A0(n4059), .A1(n7681), .B0(n6751), .B1(n4048), .Y(n5074) );
  OAI22XL U2494 ( .A0(n4061), .A1(n7809), .B0(n6751), .B1(n4072), .Y(n5202) );
  OAI22XL U2495 ( .A0(n4085), .A1(n7937), .B0(n6751), .B1(n4078), .Y(n5330) );
  OAI22XL U2496 ( .A0(n4097), .A1(n8065), .B0(n6751), .B1(n4090), .Y(n5458) );
  OAI22XL U2497 ( .A0(n4111), .A1(n8193), .B0(n6751), .B1(n4104), .Y(n5586) );
  OAI22XL U2498 ( .A0(n4185), .A1(n7297), .B0(n6751), .B1(n4179), .Y(n4690) );
  OAI22XL U2499 ( .A0(n4043), .A1(n7554), .B0(n6752), .B1(n4034), .Y(n4947) );
  OAI22XL U2500 ( .A0(n4058), .A1(n7682), .B0(n6752), .B1(n4048), .Y(n5075) );
  OAI22XL U2501 ( .A0(n4061), .A1(n7810), .B0(n6752), .B1(n4072), .Y(n5203) );
  OAI22XL U2502 ( .A0(n4085), .A1(n7938), .B0(n6752), .B1(n4078), .Y(n5331) );
  OAI22XL U2503 ( .A0(n4097), .A1(n8066), .B0(n6752), .B1(n4090), .Y(n5459) );
  OAI22XL U2504 ( .A0(n4111), .A1(n8194), .B0(n6752), .B1(n4104), .Y(n5587) );
  OAI22XL U2505 ( .A0(n4185), .A1(n7298), .B0(n6752), .B1(n4179), .Y(n4691) );
  OAI22XL U2506 ( .A0(n4043), .A1(n7555), .B0(n6753), .B1(n4034), .Y(n4948) );
  OAI22XL U2507 ( .A0(n4055), .A1(n7683), .B0(n6753), .B1(n4048), .Y(n5076) );
  OAI22XL U2508 ( .A0(n4062), .A1(n7811), .B0(n6753), .B1(n4072), .Y(n5204) );
  OAI22XL U2509 ( .A0(n4085), .A1(n7939), .B0(n6753), .B1(n4078), .Y(n5332) );
  OAI22XL U2510 ( .A0(n4097), .A1(n8067), .B0(n6753), .B1(n4090), .Y(n5460) );
  OAI22XL U2511 ( .A0(n4111), .A1(n8195), .B0(n6753), .B1(n4104), .Y(n5588) );
  OAI22XL U2512 ( .A0(n4185), .A1(n7299), .B0(n6753), .B1(n4179), .Y(n4692) );
  OAI22XL U2513 ( .A0(n4043), .A1(n7556), .B0(n6754), .B1(n4034), .Y(n4949) );
  OAI22XL U2514 ( .A0(n4053), .A1(n7684), .B0(n6754), .B1(n4048), .Y(n5077) );
  OAI22XL U2515 ( .A0(n4062), .A1(n7812), .B0(n6754), .B1(n4072), .Y(n5205) );
  OAI22XL U2516 ( .A0(n4085), .A1(n7940), .B0(n6754), .B1(n4078), .Y(n5333) );
  OAI22XL U2517 ( .A0(n4097), .A1(n8068), .B0(n6754), .B1(n4090), .Y(n5461) );
  OAI22XL U2518 ( .A0(n4111), .A1(n8196), .B0(n6754), .B1(n4104), .Y(n5589) );
  OAI22XL U2519 ( .A0(n4185), .A1(n7300), .B0(n6754), .B1(n4179), .Y(n4693) );
  OAI22XL U2520 ( .A0(n4043), .A1(n7557), .B0(n6755), .B1(n4034), .Y(n4950) );
  OAI22XL U2521 ( .A0(n4055), .A1(n7685), .B0(n6755), .B1(n4048), .Y(n5078) );
  OAI22XL U2522 ( .A0(n4062), .A1(n7813), .B0(n6755), .B1(n4072), .Y(n5206) );
  OAI22XL U2523 ( .A0(n4083), .A1(n7941), .B0(n6755), .B1(n4078), .Y(n5334) );
  OAI22XL U2524 ( .A0(n4097), .A1(n8069), .B0(n6755), .B1(n4090), .Y(n5462) );
  OAI22XL U2525 ( .A0(n4111), .A1(n8197), .B0(n6755), .B1(n4104), .Y(n5590) );
  OAI22XL U2526 ( .A0(n4186), .A1(n7301), .B0(n6755), .B1(n4180), .Y(n4694) );
  OAI22XL U2527 ( .A0(n4043), .A1(n7558), .B0(n6756), .B1(n4034), .Y(n4951) );
  OAI22XL U2528 ( .A0(n4054), .A1(n7686), .B0(n6756), .B1(n4048), .Y(n5079) );
  OAI22XL U2529 ( .A0(n4062), .A1(n7814), .B0(n6756), .B1(n4072), .Y(n5207) );
  OAI22XL U2530 ( .A0(n4082), .A1(n7942), .B0(n6756), .B1(n4078), .Y(n5335) );
  OAI22XL U2531 ( .A0(n4097), .A1(n8070), .B0(n6756), .B1(n4090), .Y(n5463) );
  OAI22XL U2532 ( .A0(n4111), .A1(n8198), .B0(n6756), .B1(n4104), .Y(n5591) );
  OAI22XL U2533 ( .A0(n4186), .A1(n7302), .B0(n6756), .B1(n4180), .Y(n4695) );
  OAI22XL U2534 ( .A0(n4043), .A1(n7559), .B0(n6757), .B1(n4034), .Y(n4952) );
  OAI22XL U2535 ( .A0(n4054), .A1(n7687), .B0(n6757), .B1(n4048), .Y(n5080) );
  OAI22XL U2536 ( .A0(n4062), .A1(n7815), .B0(n6757), .B1(n4072), .Y(n5208) );
  OAI22XL U2537 ( .A0(n4085), .A1(n7943), .B0(n6757), .B1(n4078), .Y(n5336) );
  OAI22XL U2538 ( .A0(n4097), .A1(n8071), .B0(n6757), .B1(n4090), .Y(n5464) );
  OAI22XL U2539 ( .A0(n4111), .A1(n8199), .B0(n6757), .B1(n4104), .Y(n5592) );
  OAI22XL U2540 ( .A0(n4186), .A1(n7303), .B0(n6757), .B1(n4180), .Y(n4696) );
  OAI22XL U2541 ( .A0(n4043), .A1(n7560), .B0(n6758), .B1(n4034), .Y(n4953) );
  OAI22XL U2542 ( .A0(n4055), .A1(n7688), .B0(n6758), .B1(n4048), .Y(n5081) );
  OAI22XL U2543 ( .A0(n4062), .A1(n7816), .B0(n6758), .B1(n4068), .Y(n5209) );
  OAI22XL U2544 ( .A0(n4083), .A1(n7944), .B0(n6758), .B1(n4078), .Y(n5337) );
  OAI22XL U2545 ( .A0(n4097), .A1(n8072), .B0(n6758), .B1(n4090), .Y(n5465) );
  OAI22XL U2546 ( .A0(n4111), .A1(n8200), .B0(n6758), .B1(n4104), .Y(n5593) );
  OAI22XL U2547 ( .A0(n4186), .A1(n7304), .B0(n6758), .B1(n4180), .Y(n4697) );
  OAI22XL U2548 ( .A0(n4043), .A1(n7561), .B0(n6759), .B1(n4034), .Y(n4954) );
  OAI22XL U2549 ( .A0(n4054), .A1(n7689), .B0(n6759), .B1(n4048), .Y(n5082) );
  OAI22XL U2550 ( .A0(n4062), .A1(n7817), .B0(n6759), .B1(n4072), .Y(n5210) );
  OAI22XL U2551 ( .A0(n4083), .A1(n7945), .B0(n6759), .B1(n4077), .Y(n5338) );
  OAI22XL U2552 ( .A0(n4097), .A1(n8073), .B0(n6759), .B1(n4090), .Y(n5466) );
  OAI22XL U2553 ( .A0(n4111), .A1(n8201), .B0(n6759), .B1(n4104), .Y(n5594) );
  OAI22XL U2554 ( .A0(n4186), .A1(n7305), .B0(n6759), .B1(n4180), .Y(n4698) );
  OAI22XL U2555 ( .A0(n4043), .A1(n7562), .B0(n6760), .B1(n4034), .Y(n4955) );
  OAI22XL U2556 ( .A0(n4057), .A1(n7690), .B0(n6760), .B1(n4048), .Y(n5083) );
  OAI22XL U2557 ( .A0(n4062), .A1(n7818), .B0(n6760), .B1(n4068), .Y(n5211) );
  OAI22XL U2558 ( .A0(n4084), .A1(n7946), .B0(n6760), .B1(n4077), .Y(n5339) );
  OAI22XL U2559 ( .A0(n4097), .A1(n8074), .B0(n6760), .B1(n4090), .Y(n5467) );
  OAI22XL U2560 ( .A0(n4111), .A1(n8202), .B0(n6760), .B1(n4104), .Y(n5595) );
  OAI22XL U2561 ( .A0(n4186), .A1(n7306), .B0(n6760), .B1(n4180), .Y(n4699) );
  OAI22XL U2562 ( .A0(n4044), .A1(n7563), .B0(n6761), .B1(n4035), .Y(n4956) );
  OAI22XL U2563 ( .A0(n4055), .A1(n7691), .B0(n6761), .B1(n4049), .Y(n5084) );
  OAI22XL U2564 ( .A0(n4062), .A1(n7819), .B0(n6761), .B1(n4072), .Y(n5212) );
  OAI22XL U2565 ( .A0(n4081), .A1(n7947), .B0(n6761), .B1(n4077), .Y(n5340) );
  OAI22XL U2566 ( .A0(n4094), .A1(n8075), .B0(n6761), .B1(n4091), .Y(n5468) );
  OAI22XL U2567 ( .A0(n4108), .A1(n8203), .B0(n6761), .B1(n4105), .Y(n5596) );
  OAI22XL U2568 ( .A0(n4186), .A1(n7307), .B0(n6761), .B1(n4180), .Y(n4700) );
  OAI22XL U2569 ( .A0(n4044), .A1(n7564), .B0(n6762), .B1(n4035), .Y(n4957) );
  OAI22XL U2570 ( .A0(n4055), .A1(n7692), .B0(n6762), .B1(n4049), .Y(n5085) );
  OAI22XL U2571 ( .A0(n4062), .A1(n7820), .B0(n6762), .B1(n4068), .Y(n5213) );
  OAI22XL U2572 ( .A0(n4085), .A1(n7948), .B0(n6762), .B1(n4077), .Y(n5341) );
  OAI22XL U2573 ( .A0(n4093), .A1(n8076), .B0(n6762), .B1(n4091), .Y(n5469) );
  OAI22XL U2574 ( .A0(n4107), .A1(n8204), .B0(n6762), .B1(n4105), .Y(n5597) );
  OAI22XL U2575 ( .A0(n4186), .A1(n7308), .B0(n6762), .B1(n4180), .Y(n4701) );
  OAI22XL U2576 ( .A0(n4044), .A1(n7565), .B0(n6763), .B1(n4035), .Y(n4958) );
  OAI22XL U2577 ( .A0(n4055), .A1(n7693), .B0(n6763), .B1(n4049), .Y(n5086) );
  OAI22XL U2578 ( .A0(n4062), .A1(n7821), .B0(n6763), .B1(n4072), .Y(n5214) );
  OAI22XL U2579 ( .A0(n4083), .A1(n7949), .B0(n6763), .B1(n4077), .Y(n5342) );
  OAI22XL U2580 ( .A0(n4099), .A1(n8077), .B0(n6763), .B1(n4091), .Y(n5470) );
  OAI22XL U2581 ( .A0(n4113), .A1(n8205), .B0(n6763), .B1(n4105), .Y(n5598) );
  OAI22XL U2582 ( .A0(n4186), .A1(n7309), .B0(n6763), .B1(n4180), .Y(n4702) );
  OAI22XL U2583 ( .A0(n4044), .A1(n7566), .B0(n6764), .B1(n4035), .Y(n4959) );
  OAI22XL U2584 ( .A0(n4055), .A1(n7694), .B0(n6764), .B1(n4049), .Y(n5087) );
  OAI22XL U2585 ( .A0(n4062), .A1(n7822), .B0(n6764), .B1(n4068), .Y(n5215) );
  OAI22XL U2586 ( .A0(n4082), .A1(n7950), .B0(n6764), .B1(n4077), .Y(n5343) );
  OAI22XL U2587 ( .A0(n4099), .A1(n8078), .B0(n6764), .B1(n4091), .Y(n5471) );
  OAI22XL U2588 ( .A0(n4113), .A1(n8206), .B0(n6764), .B1(n4105), .Y(n5599) );
  OAI22XL U2589 ( .A0(n4186), .A1(n7310), .B0(n6764), .B1(n4180), .Y(n4703) );
  OAI22XL U2590 ( .A0(n4044), .A1(n7567), .B0(n6765), .B1(n4035), .Y(n4960) );
  OAI22XL U2591 ( .A0(n4055), .A1(n7695), .B0(n6765), .B1(n4049), .Y(n5088) );
  OAI22XL U2592 ( .A0(n4063), .A1(n7823), .B0(n6765), .B1(n4067), .Y(n5216) );
  OAI22XL U2593 ( .A0(n4084), .A1(n7951), .B0(n6765), .B1(n4077), .Y(n5344) );
  OAI22XL U2594 ( .A0(n4099), .A1(n8079), .B0(n6765), .B1(n4091), .Y(n5472) );
  OAI22XL U2595 ( .A0(n4113), .A1(n8207), .B0(n6765), .B1(n4105), .Y(n5600) );
  OAI22XL U2596 ( .A0(n4186), .A1(n7311), .B0(n6765), .B1(n4180), .Y(n4704) );
  OAI22XL U2597 ( .A0(n4044), .A1(n7568), .B0(n6766), .B1(n4035), .Y(n4961) );
  OAI22XL U2598 ( .A0(n4055), .A1(n7696), .B0(n6766), .B1(n4049), .Y(n5089) );
  OAI22XL U2599 ( .A0(n4063), .A1(n7824), .B0(n6766), .B1(n4067), .Y(n5217) );
  OAI22XL U2600 ( .A0(n4084), .A1(n7952), .B0(n6766), .B1(n4077), .Y(n5345) );
  OAI22XL U2601 ( .A0(n4099), .A1(n8080), .B0(n6766), .B1(n4091), .Y(n5473) );
  OAI22XL U2602 ( .A0(n4113), .A1(n8208), .B0(n6766), .B1(n4105), .Y(n5601) );
  OAI22XL U2603 ( .A0(n4186), .A1(n7312), .B0(n6766), .B1(n4180), .Y(n4705) );
  OAI22XL U2604 ( .A0(n4044), .A1(n7569), .B0(n6767), .B1(n4035), .Y(n4962) );
  OAI22XL U2605 ( .A0(n4055), .A1(n7697), .B0(n6767), .B1(n4049), .Y(n5090) );
  OAI22XL U2606 ( .A0(n4063), .A1(n7825), .B0(n6767), .B1(n4070), .Y(n5218) );
  OAI22XL U2607 ( .A0(n4081), .A1(n7953), .B0(n6767), .B1(n4077), .Y(n5346) );
  OAI22XL U2608 ( .A0(n4095), .A1(n8081), .B0(n6767), .B1(n4091), .Y(n5474) );
  OAI22XL U2609 ( .A0(n4109), .A1(n8209), .B0(n6767), .B1(n4105), .Y(n5602) );
  OAI22XL U2610 ( .A0(n4187), .A1(n7313), .B0(n6767), .B1(n4184), .Y(n4706) );
  OAI22XL U2611 ( .A0(n4044), .A1(n7570), .B0(n6768), .B1(n4035), .Y(n4963) );
  OAI22XL U2612 ( .A0(n4055), .A1(n7698), .B0(n6768), .B1(n4049), .Y(n5091) );
  OAI22XL U2613 ( .A0(n4063), .A1(n7826), .B0(n6768), .B1(n4071), .Y(n5219) );
  OAI22XL U2614 ( .A0(n4081), .A1(n7954), .B0(n6768), .B1(n4077), .Y(n5347) );
  OAI22XL U2615 ( .A0(n4098), .A1(n8082), .B0(n6768), .B1(n4091), .Y(n5475) );
  OAI22XL U2616 ( .A0(n4112), .A1(n8210), .B0(n6768), .B1(n4105), .Y(n5603) );
  OAI22XL U2617 ( .A0(n4187), .A1(n7314), .B0(n6768), .B1(n4184), .Y(n4707) );
  OAI22XL U2618 ( .A0(n4044), .A1(n7571), .B0(n6769), .B1(n4035), .Y(n4964) );
  OAI22XL U2619 ( .A0(n4055), .A1(n7699), .B0(n6769), .B1(n4049), .Y(n5092) );
  OAI22XL U2620 ( .A0(n4063), .A1(n7827), .B0(n6769), .B1(n4067), .Y(n5220) );
  OAI22XL U2621 ( .A0(n4081), .A1(n7955), .B0(n6769), .B1(n4077), .Y(n5348) );
  OAI22XL U2622 ( .A0(n4096), .A1(n8083), .B0(n6769), .B1(n4091), .Y(n5476) );
  OAI22XL U2623 ( .A0(n4110), .A1(n8211), .B0(n6769), .B1(n4105), .Y(n5604) );
  OAI22XL U2624 ( .A0(n4187), .A1(n7315), .B0(n6769), .B1(n4184), .Y(n4708) );
  OAI22XL U2625 ( .A0(n4044), .A1(n7572), .B0(n6770), .B1(n4035), .Y(n4965) );
  OAI22XL U2626 ( .A0(n4055), .A1(n7700), .B0(n6770), .B1(n4049), .Y(n5093) );
  OAI22XL U2627 ( .A0(n4063), .A1(n7828), .B0(n6770), .B1(n4071), .Y(n5221) );
  OAI22XL U2628 ( .A0(n4081), .A1(n7956), .B0(n6770), .B1(n4077), .Y(n5349) );
  OAI22XL U2629 ( .A0(n4097), .A1(n8084), .B0(n6770), .B1(n4091), .Y(n5477) );
  OAI22XL U2630 ( .A0(n4111), .A1(n8212), .B0(n6770), .B1(n4105), .Y(n5605) );
  OAI22XL U2631 ( .A0(n4187), .A1(n7316), .B0(n6770), .B1(n4184), .Y(n4709) );
  OAI22XL U2632 ( .A0(n4044), .A1(n7573), .B0(n6771), .B1(n4035), .Y(n4966) );
  OAI22XL U2633 ( .A0(n4055), .A1(n7701), .B0(n6771), .B1(n4049), .Y(n5094) );
  OAI22XL U2634 ( .A0(n4063), .A1(n7829), .B0(n6771), .B1(n4071), .Y(n5222) );
  OAI22XL U2635 ( .A0(n6715), .A1(n7957), .B0(n6771), .B1(n4076), .Y(n5350) );
  OAI22XL U2636 ( .A0(n4094), .A1(n8085), .B0(n6771), .B1(n4091), .Y(n5478) );
  OAI22XL U2637 ( .A0(n4108), .A1(n8213), .B0(n6771), .B1(n4105), .Y(n5606) );
  OAI22XL U2638 ( .A0(n4187), .A1(n7317), .B0(n6771), .B1(n4184), .Y(n4710) );
  OAI22XL U2639 ( .A0(n4044), .A1(n7574), .B0(n6772), .B1(n4035), .Y(n4967) );
  OAI22XL U2640 ( .A0(n4055), .A1(n7702), .B0(n6772), .B1(n4049), .Y(n5095) );
  OAI22XL U2641 ( .A0(n4063), .A1(n7830), .B0(n6772), .B1(n4071), .Y(n5223) );
  OAI22XL U2642 ( .A0(n6715), .A1(n7958), .B0(n6772), .B1(n4076), .Y(n5351) );
  OAI22XL U2643 ( .A0(n4093), .A1(n8086), .B0(n6772), .B1(n4091), .Y(n5479) );
  OAI22XL U2644 ( .A0(n4107), .A1(n8214), .B0(n6772), .B1(n4105), .Y(n5607) );
  OAI22XL U2645 ( .A0(n4187), .A1(n7318), .B0(n6772), .B1(n4184), .Y(n4711) );
  OAI22XL U2646 ( .A0(n4042), .A1(n7575), .B0(n6773), .B1(n4036), .Y(n4968) );
  OAI22XL U2647 ( .A0(n6712), .A1(n7703), .B0(n6773), .B1(n4049), .Y(n5096) );
  OAI22XL U2648 ( .A0(n4063), .A1(n7831), .B0(n6773), .B1(n4071), .Y(n5224) );
  OAI22XL U2649 ( .A0(n6715), .A1(n7959), .B0(n6773), .B1(n4076), .Y(n5352) );
  OAI22XL U2650 ( .A0(n4098), .A1(n8087), .B0(n6773), .B1(n4091), .Y(n5480) );
  OAI22XL U2651 ( .A0(n4112), .A1(n8215), .B0(n6773), .B1(n4105), .Y(n5608) );
  OAI22XL U2652 ( .A0(n4187), .A1(n7319), .B0(n6773), .B1(n4184), .Y(n4712) );
  OAI22XL U2653 ( .A0(n4040), .A1(n7576), .B0(n6774), .B1(n4036), .Y(n4969) );
  OAI22XL U2654 ( .A0(n6712), .A1(n7704), .B0(n6774), .B1(n4052), .Y(n5097) );
  OAI22XL U2655 ( .A0(n4063), .A1(n7832), .B0(n6774), .B1(n4071), .Y(n5225) );
  OAI22XL U2656 ( .A0(n6715), .A1(n7960), .B0(n6774), .B1(n4076), .Y(n5353) );
  OAI22XL U2657 ( .A0(n4098), .A1(n8088), .B0(n6774), .B1(n4088), .Y(n5481) );
  OAI22XL U2658 ( .A0(n4112), .A1(n8216), .B0(n6774), .B1(n4102), .Y(n5609) );
  OAI22XL U2659 ( .A0(n4187), .A1(n7320), .B0(n6774), .B1(n4182), .Y(n4713) );
  OAI22XL U2660 ( .A0(n4044), .A1(n7577), .B0(n6775), .B1(n4036), .Y(n4970) );
  OAI22XL U2661 ( .A0(n6712), .A1(n7705), .B0(n6775), .B1(n4052), .Y(n5098) );
  OAI22XL U2662 ( .A0(n4063), .A1(n7833), .B0(n6775), .B1(n4071), .Y(n5226) );
  OAI22XL U2663 ( .A0(n6715), .A1(n7961), .B0(n6775), .B1(n4076), .Y(n5354) );
  OAI22XL U2664 ( .A0(n4098), .A1(n8089), .B0(n6775), .B1(n4087), .Y(n5482) );
  OAI22XL U2665 ( .A0(n4112), .A1(n8217), .B0(n6775), .B1(n4101), .Y(n5610) );
  OAI22XL U2666 ( .A0(n4187), .A1(n7321), .B0(n6775), .B1(n4182), .Y(n4714) );
  OAI22XL U2667 ( .A0(n4044), .A1(n7578), .B0(n6776), .B1(n4036), .Y(n4971) );
  OAI22XL U2668 ( .A0(n6712), .A1(n7706), .B0(n6776), .B1(n4052), .Y(n5099) );
  OAI22XL U2669 ( .A0(n4063), .A1(n7834), .B0(n6776), .B1(n4071), .Y(n5227) );
  OAI22XL U2670 ( .A0(n4081), .A1(n7962), .B0(n6776), .B1(n4076), .Y(n5355) );
  OAI22XL U2671 ( .A0(n4098), .A1(n8090), .B0(n6776), .B1(n4087), .Y(n5483) );
  OAI22XL U2672 ( .A0(n4112), .A1(n8218), .B0(n6776), .B1(n4101), .Y(n5611) );
  OAI22XL U2673 ( .A0(n4187), .A1(n7322), .B0(n6776), .B1(n4182), .Y(n4715) );
  OAI22XL U2674 ( .A0(n4044), .A1(n7579), .B0(n6777), .B1(n4036), .Y(n4972) );
  OAI22XL U2675 ( .A0(n6712), .A1(n7707), .B0(n6777), .B1(n4052), .Y(n5100) );
  OAI22XL U2676 ( .A0(n4064), .A1(n7835), .B0(n6777), .B1(n4071), .Y(n5228) );
  OAI22XL U2677 ( .A0(n4081), .A1(n7963), .B0(n6777), .B1(n4076), .Y(n5356) );
  OAI22XL U2678 ( .A0(n4098), .A1(n8091), .B0(n6777), .B1(n4087), .Y(n5484) );
  OAI22XL U2679 ( .A0(n4112), .A1(n8219), .B0(n6777), .B1(n4101), .Y(n5612) );
  OAI22XL U2680 ( .A0(n4187), .A1(n7323), .B0(n6777), .B1(n4179), .Y(n4716) );
  OAI22XL U2681 ( .A0(n4039), .A1(n7580), .B0(n6778), .B1(n4036), .Y(n4973) );
  OAI22XL U2682 ( .A0(n4053), .A1(n7708), .B0(n6778), .B1(n4052), .Y(n5101) );
  OAI22XL U2683 ( .A0(n4064), .A1(n7836), .B0(n6778), .B1(n4071), .Y(n5229) );
  OAI22XL U2684 ( .A0(n4081), .A1(n7964), .B0(n6778), .B1(n4076), .Y(n5357) );
  OAI22XL U2685 ( .A0(n4098), .A1(n8092), .B0(n6778), .B1(n4087), .Y(n5485) );
  OAI22XL U2686 ( .A0(n4112), .A1(n8220), .B0(n6778), .B1(n4101), .Y(n5613) );
  OAI22XL U2687 ( .A0(n4187), .A1(n7324), .B0(n6778), .B1(n4180), .Y(n4717) );
  OAI22XL U2688 ( .A0(n4039), .A1(n7581), .B0(n6779), .B1(n4036), .Y(n4974) );
  OAI22XL U2689 ( .A0(n4053), .A1(n7709), .B0(n6779), .B1(n4052), .Y(n5102) );
  OAI22XL U2690 ( .A0(n4064), .A1(n7837), .B0(n6779), .B1(n4071), .Y(n5230) );
  OAI22XL U2691 ( .A0(n4081), .A1(n7965), .B0(n6779), .B1(n4076), .Y(n5358) );
  OAI22XL U2692 ( .A0(n4098), .A1(n8093), .B0(n6779), .B1(n4087), .Y(n5486) );
  OAI22XL U2693 ( .A0(n4112), .A1(n8221), .B0(n6779), .B1(n4101), .Y(n5614) );
  OAI22XL U2694 ( .A0(n4187), .A1(n7325), .B0(n6779), .B1(n4181), .Y(n4718) );
  OAI22XL U2695 ( .A0(n4039), .A1(n7582), .B0(n6780), .B1(n4036), .Y(n4975) );
  OAI22XL U2696 ( .A0(n4053), .A1(n7710), .B0(n6780), .B1(n4052), .Y(n5103) );
  OAI22XL U2697 ( .A0(n4064), .A1(n7838), .B0(n6780), .B1(n4071), .Y(n5231) );
  OAI22XL U2698 ( .A0(n4085), .A1(n7966), .B0(n6780), .B1(n4076), .Y(n5359) );
  OAI22XL U2699 ( .A0(n4098), .A1(n8094), .B0(n6780), .B1(n4089), .Y(n5487) );
  OAI22XL U2700 ( .A0(n4112), .A1(n8222), .B0(n6780), .B1(n4103), .Y(n5615) );
  OAI22XL U2701 ( .A0(n4186), .A1(n7326), .B0(n6780), .B1(n4181), .Y(n4719) );
  OAI22XL U2702 ( .A0(n4039), .A1(n7583), .B0(n6781), .B1(n4036), .Y(n4976) );
  OAI22XL U2703 ( .A0(n4053), .A1(n7711), .B0(n6781), .B1(n4052), .Y(n5104) );
  OAI22XL U2704 ( .A0(n4064), .A1(n7839), .B0(n6781), .B1(n4071), .Y(n5232) );
  OAI22XL U2705 ( .A0(n4083), .A1(n7967), .B0(n6781), .B1(n4076), .Y(n5360) );
  OAI22XL U2706 ( .A0(n4098), .A1(n8095), .B0(n6781), .B1(n4090), .Y(n5488) );
  OAI22XL U2707 ( .A0(n4112), .A1(n8223), .B0(n6781), .B1(n4104), .Y(n5616) );
  OAI22XL U2708 ( .A0(n4189), .A1(n7327), .B0(n6781), .B1(n4181), .Y(n4720) );
  OAI22XL U2709 ( .A0(n6711), .A1(n7584), .B0(n6782), .B1(n4036), .Y(n4977) );
  OAI22XL U2710 ( .A0(n4053), .A1(n7712), .B0(n6782), .B1(n4052), .Y(n5105) );
  OAI22XL U2711 ( .A0(n4064), .A1(n7840), .B0(n6782), .B1(n4070), .Y(n5233) );
  OAI22XL U2712 ( .A0(n4084), .A1(n7968), .B0(n6782), .B1(n4076), .Y(n5361) );
  OAI22XL U2713 ( .A0(n4098), .A1(n8096), .B0(n6782), .B1(n4091), .Y(n5489) );
  OAI22XL U2714 ( .A0(n4112), .A1(n8224), .B0(n6782), .B1(n4105), .Y(n5617) );
  OAI22XL U2715 ( .A0(n4187), .A1(n7328), .B0(n6782), .B1(n4181), .Y(n4721) );
  OAI22XL U2716 ( .A0(n6711), .A1(n7585), .B0(n6783), .B1(n4036), .Y(n4978) );
  OAI22XL U2717 ( .A0(n4053), .A1(n7713), .B0(n6783), .B1(n4052), .Y(n5106) );
  OAI22XL U2718 ( .A0(n4064), .A1(n7841), .B0(n6783), .B1(n4070), .Y(n5234) );
  OAI22XL U2719 ( .A0(n4082), .A1(n7969), .B0(n6783), .B1(n4076), .Y(n5362) );
  OAI22XL U2720 ( .A0(n4098), .A1(n8097), .B0(n6783), .B1(n4088), .Y(n5490) );
  OAI22XL U2721 ( .A0(n4112), .A1(n8225), .B0(n6783), .B1(n4102), .Y(n5618) );
  OAI22XL U2722 ( .A0(n4187), .A1(n7329), .B0(n6783), .B1(n4181), .Y(n4722) );
  OAI22XL U2723 ( .A0(n6711), .A1(n7586), .B0(n6784), .B1(n4036), .Y(n4979) );
  OAI22XL U2724 ( .A0(n4053), .A1(n7714), .B0(n6784), .B1(n4052), .Y(n5107) );
  OAI22XL U2725 ( .A0(n4064), .A1(n7842), .B0(n6784), .B1(n4070), .Y(n5235) );
  OAI22XL U2726 ( .A0(n4085), .A1(n7970), .B0(n6784), .B1(n4076), .Y(n5363) );
  OAI22XL U2727 ( .A0(n4098), .A1(n8098), .B0(n6784), .B1(n4089), .Y(n5491) );
  OAI22XL U2728 ( .A0(n4112), .A1(n8226), .B0(n6784), .B1(n4103), .Y(n5619) );
  OAI22XL U2729 ( .A0(n4186), .A1(n7330), .B0(n6784), .B1(n4181), .Y(n4723) );
  OAI22XL U2730 ( .A0(n4039), .A1(n7587), .B0(n6785), .B1(n4037), .Y(n4980) );
  OAI22XL U2731 ( .A0(n4056), .A1(n7715), .B0(n6785), .B1(n4050), .Y(n5108) );
  OAI22XL U2732 ( .A0(n4064), .A1(n7843), .B0(n6785), .B1(n4070), .Y(n5236) );
  OAI22XL U2733 ( .A0(n4083), .A1(n7971), .B0(n6785), .B1(n4078), .Y(n5364) );
  OAI22XL U2734 ( .A0(n4095), .A1(n8099), .B0(n6785), .B1(n4088), .Y(n5492) );
  OAI22XL U2735 ( .A0(n4109), .A1(n8227), .B0(n6785), .B1(n4102), .Y(n5620) );
  OAI22XL U2736 ( .A0(n4189), .A1(n7331), .B0(n6785), .B1(n4181), .Y(n4724) );
  OAI22XL U2737 ( .A0(n4039), .A1(n7588), .B0(n6786), .B1(n4037), .Y(n4981) );
  OAI22XL U2738 ( .A0(n4056), .A1(n7716), .B0(n6786), .B1(n4050), .Y(n5109) );
  OAI22XL U2739 ( .A0(n4064), .A1(n7844), .B0(n6786), .B1(n4070), .Y(n5237) );
  OAI22XL U2740 ( .A0(n4084), .A1(n7972), .B0(n6786), .B1(n4076), .Y(n5365) );
  OAI22XL U2741 ( .A0(n4099), .A1(n8100), .B0(n6786), .B1(n4091), .Y(n5493) );
  OAI22XL U2742 ( .A0(n4113), .A1(n8228), .B0(n6786), .B1(n4105), .Y(n5621) );
  OAI22XL U2743 ( .A0(n4186), .A1(n7332), .B0(n6786), .B1(n4181), .Y(n4725) );
  OAI22XL U2744 ( .A0(n4039), .A1(n7589), .B0(n6787), .B1(n4037), .Y(n4982) );
  OAI22XL U2745 ( .A0(n4056), .A1(n7717), .B0(n6787), .B1(n4050), .Y(n5110) );
  OAI22XL U2746 ( .A0(n4064), .A1(n7845), .B0(n6787), .B1(n4070), .Y(n5238) );
  OAI22XL U2747 ( .A0(n4082), .A1(n7973), .B0(n6787), .B1(n4078), .Y(n5366) );
  OAI22XL U2748 ( .A0(n4098), .A1(n8101), .B0(n6787), .B1(n4090), .Y(n5494) );
  OAI22XL U2749 ( .A0(n4112), .A1(n8229), .B0(n6787), .B1(n4104), .Y(n5622) );
  OAI22XL U2750 ( .A0(n4187), .A1(n7333), .B0(n6787), .B1(n4181), .Y(n4726) );
  OAI22XL U2751 ( .A0(n4039), .A1(n7590), .B0(n6788), .B1(n4037), .Y(n4983) );
  OAI22XL U2752 ( .A0(n4056), .A1(n7718), .B0(n6788), .B1(n4050), .Y(n5111) );
  OAI22XL U2753 ( .A0(n4064), .A1(n7846), .B0(n6788), .B1(n4070), .Y(n5239) );
  OAI22XL U2754 ( .A0(n4084), .A1(n7974), .B0(n6788), .B1(n4079), .Y(n5367) );
  OAI22XL U2755 ( .A0(n4096), .A1(n8102), .B0(n6788), .B1(n4089), .Y(n5495) );
  OAI22XL U2756 ( .A0(n4110), .A1(n8230), .B0(n6788), .B1(n4103), .Y(n5623) );
  OAI22XL U2757 ( .A0(n4186), .A1(n7334), .B0(n6788), .B1(n4181), .Y(n4727) );
  OAI22XL U2758 ( .A0(n4039), .A1(n7591), .B0(n6789), .B1(n4037), .Y(n4984) );
  OAI22XL U2759 ( .A0(n4056), .A1(n7719), .B0(n6789), .B1(n4050), .Y(n5112) );
  OAI22XL U2760 ( .A0(n4065), .A1(n7847), .B0(n6789), .B1(n4070), .Y(n5240) );
  OAI22XL U2761 ( .A0(n4085), .A1(n7975), .B0(n6789), .B1(n4076), .Y(n5368) );
  OAI22XL U2762 ( .A0(n4097), .A1(n8103), .B0(n6789), .B1(n4090), .Y(n5496) );
  OAI22XL U2763 ( .A0(n4111), .A1(n8231), .B0(n6789), .B1(n4104), .Y(n5624) );
  OAI22XL U2764 ( .A0(n4189), .A1(n7335), .B0(n6789), .B1(n4181), .Y(n4728) );
  OAI22XL U2765 ( .A0(n4039), .A1(n7509), .B0(n6868), .B1(n4038), .Y(n4902) );
  OAI22XL U2766 ( .A0(n4053), .A1(n7637), .B0(n6868), .B1(n4052), .Y(n5030) );
  OAI22XL U2767 ( .A0(n4062), .A1(n7765), .B0(n6868), .B1(n4073), .Y(n5158) );
  OAI22XL U2768 ( .A0(n4082), .A1(n7893), .B0(n6868), .B1(n4078), .Y(n5286) );
  OAI22XL U2769 ( .A0(n4093), .A1(n8021), .B0(n6868), .B1(n4086), .Y(n5414) );
  OAI22XL U2770 ( .A0(n4107), .A1(n8149), .B0(n6868), .B1(n4100), .Y(n5542) );
  OAI22XL U2771 ( .A0(n4185), .A1(n7253), .B0(n6868), .B1(n4184), .Y(n4646) );
  OAI22XL U2772 ( .A0(n4043), .A1(n7510), .B0(n6869), .B1(n4033), .Y(n4903) );
  OAI22XL U2773 ( .A0(n4057), .A1(n7638), .B0(n6869), .B1(n4048), .Y(n5031) );
  OAI22XL U2774 ( .A0(n4063), .A1(n7766), .B0(n6869), .B1(n4073), .Y(n5159) );
  OAI22XL U2775 ( .A0(n4082), .A1(n7894), .B0(n6869), .B1(n4074), .Y(n5287) );
  OAI22XL U2776 ( .A0(n4093), .A1(n8022), .B0(n6869), .B1(n4086), .Y(n5415) );
  OAI22XL U2777 ( .A0(n4107), .A1(n8150), .B0(n6869), .B1(n4100), .Y(n5543) );
  OAI22XL U2778 ( .A0(n4191), .A1(n7254), .B0(n6869), .B1(n4184), .Y(n4647) );
  OAI22XL U2779 ( .A0(n4041), .A1(n7511), .B0(n6870), .B1(n4034), .Y(n4904) );
  OAI22XL U2780 ( .A0(n4059), .A1(n7639), .B0(n6870), .B1(n4047), .Y(n5032) );
  OAI22XL U2781 ( .A0(n4064), .A1(n7767), .B0(n6870), .B1(n4073), .Y(n5160) );
  OAI22XL U2782 ( .A0(n4082), .A1(n7895), .B0(n6870), .B1(n4080), .Y(n5288) );
  OAI22XL U2783 ( .A0(n4093), .A1(n8023), .B0(n6870), .B1(n4086), .Y(n5416) );
  OAI22XL U2784 ( .A0(n4107), .A1(n8151), .B0(n6870), .B1(n4100), .Y(n5544) );
  OAI22XL U2785 ( .A0(n4189), .A1(n7255), .B0(n6870), .B1(n4184), .Y(n4648) );
  OAI22XL U2786 ( .A0(n4039), .A1(n7512), .B0(n6871), .B1(n4036), .Y(n4905) );
  OAI22XL U2787 ( .A0(n4053), .A1(n7640), .B0(n6871), .B1(n4046), .Y(n5033) );
  OAI22XL U2788 ( .A0(n4065), .A1(n7768), .B0(n6871), .B1(n4073), .Y(n5161) );
  OAI22XL U2789 ( .A0(n4082), .A1(n7896), .B0(n6871), .B1(n4074), .Y(n5289) );
  OAI22XL U2790 ( .A0(n4093), .A1(n8024), .B0(n6871), .B1(n4086), .Y(n5417) );
  OAI22XL U2791 ( .A0(n4107), .A1(n8152), .B0(n6871), .B1(n4100), .Y(n5545) );
  OAI22XL U2792 ( .A0(n4191), .A1(n7256), .B0(n6871), .B1(n4184), .Y(n4649) );
  OAI22XL U2793 ( .A0(n4039), .A1(n7513), .B0(n6872), .B1(n4032), .Y(n4906) );
  OAI22XL U2794 ( .A0(n4056), .A1(n7641), .B0(n6872), .B1(n4049), .Y(n5034) );
  OAI22XL U2795 ( .A0(n4061), .A1(n7769), .B0(n6872), .B1(n4073), .Y(n5162) );
  OAI22XL U2796 ( .A0(n4082), .A1(n7897), .B0(n6872), .B1(n4080), .Y(n5290) );
  OAI22XL U2797 ( .A0(n4093), .A1(n8025), .B0(n6872), .B1(n4086), .Y(n5418) );
  OAI22XL U2798 ( .A0(n4107), .A1(n8153), .B0(n6872), .B1(n4100), .Y(n5546) );
  OAI22XL U2799 ( .A0(n4188), .A1(n7257), .B0(n6872), .B1(n4178), .Y(n4650) );
  OAI22XL U2800 ( .A0(n4042), .A1(n7514), .B0(n6873), .B1(n4037), .Y(n4907) );
  OAI22XL U2801 ( .A0(n4059), .A1(n7642), .B0(n6873), .B1(n4051), .Y(n5035) );
  OAI22XL U2802 ( .A0(n4062), .A1(n7770), .B0(n6873), .B1(n4073), .Y(n5163) );
  OAI22XL U2803 ( .A0(n4082), .A1(n7898), .B0(n6873), .B1(n4074), .Y(n5291) );
  OAI22XL U2804 ( .A0(n4093), .A1(n8026), .B0(n6873), .B1(n4086), .Y(n5419) );
  OAI22XL U2805 ( .A0(n4107), .A1(n8154), .B0(n6873), .B1(n4100), .Y(n5547) );
  OAI22XL U2806 ( .A0(n4188), .A1(n7258), .B0(n6873), .B1(n4184), .Y(n4651) );
  OAI22XL U2807 ( .A0(n4040), .A1(n7515), .B0(n6874), .B1(n4032), .Y(n4908) );
  OAI22XL U2808 ( .A0(n4059), .A1(n7643), .B0(n6874), .B1(n4051), .Y(n5036) );
  OAI22XL U2809 ( .A0(n6713), .A1(n7771), .B0(n6874), .B1(n4073), .Y(n5164) );
  OAI22XL U2810 ( .A0(n4082), .A1(n7899), .B0(n6874), .B1(n4080), .Y(n5292) );
  OAI22XL U2811 ( .A0(n4094), .A1(n8027), .B0(n6874), .B1(n4087), .Y(n5420) );
  OAI22XL U2812 ( .A0(n4108), .A1(n8155), .B0(n6874), .B1(n4101), .Y(n5548) );
  OAI22XL U2813 ( .A0(n4185), .A1(n7259), .B0(n6874), .B1(n4183), .Y(n4652) );
  OAI22XL U2814 ( .A0(n4040), .A1(n7516), .B0(n6875), .B1(n4032), .Y(n4909) );
  OAI22XL U2815 ( .A0(n4057), .A1(n7644), .B0(n6875), .B1(n4046), .Y(n5037) );
  OAI22XL U2816 ( .A0(n6713), .A1(n7772), .B0(n6875), .B1(n4073), .Y(n5165) );
  OAI22XL U2817 ( .A0(n4082), .A1(n7900), .B0(n6875), .B1(n4074), .Y(n5293) );
  OAI22XL U2818 ( .A0(n4094), .A1(n8028), .B0(n6875), .B1(n4087), .Y(n5421) );
  OAI22XL U2819 ( .A0(n4108), .A1(n8156), .B0(n6875), .B1(n4101), .Y(n5549) );
  OAI22XL U2820 ( .A0(n4188), .A1(n7260), .B0(n6875), .B1(n4183), .Y(n4653) );
  OAI22XL U2821 ( .A0(n4040), .A1(n7517), .B0(n6876), .B1(n4037), .Y(n4910) );
  OAI22XL U2822 ( .A0(n4059), .A1(n7645), .B0(n6876), .B1(n4050), .Y(n5038) );
  OAI22XL U2823 ( .A0(n6713), .A1(n7773), .B0(n6876), .B1(n4069), .Y(n5166) );
  OAI22XL U2824 ( .A0(n4082), .A1(n7901), .B0(n6876), .B1(n4080), .Y(n5294) );
  OAI22XL U2825 ( .A0(n4094), .A1(n8029), .B0(n6876), .B1(n4087), .Y(n5422) );
  OAI22XL U2826 ( .A0(n4108), .A1(n8157), .B0(n6876), .B1(n4101), .Y(n5550) );
  OAI22XL U2827 ( .A0(n4190), .A1(n7261), .B0(n6876), .B1(n4182), .Y(n4654) );
  OAI22XL U2828 ( .A0(n4040), .A1(n7518), .B0(n6877), .B1(n4035), .Y(n4911) );
  OAI22XL U2829 ( .A0(n4059), .A1(n7646), .B0(n6877), .B1(n4049), .Y(n5039) );
  OAI22XL U2830 ( .A0(n6713), .A1(n7774), .B0(n6877), .B1(n4067), .Y(n5167) );
  OAI22XL U2831 ( .A0(n4082), .A1(n7902), .B0(n6877), .B1(n4074), .Y(n5295) );
  OAI22XL U2832 ( .A0(n4094), .A1(n8030), .B0(n6877), .B1(n4087), .Y(n5423) );
  OAI22XL U2833 ( .A0(n4108), .A1(n8158), .B0(n6877), .B1(n4101), .Y(n5551) );
  OAI22XL U2834 ( .A0(n4188), .A1(n7262), .B0(n6877), .B1(n4183), .Y(n4655) );
  OAI22XL U2835 ( .A0(n4040), .A1(n7519), .B0(n6878), .B1(n4038), .Y(n4912) );
  OAI22XL U2836 ( .A0(n4055), .A1(n7647), .B0(n6878), .B1(n4052), .Y(n5040) );
  OAI22XL U2837 ( .A0(n6713), .A1(n7775), .B0(n6878), .B1(n4070), .Y(n5168) );
  OAI22XL U2838 ( .A0(n4082), .A1(n7903), .B0(n6878), .B1(n4080), .Y(n5296) );
  OAI22XL U2839 ( .A0(n4094), .A1(n8031), .B0(n6878), .B1(n4087), .Y(n5424) );
  OAI22XL U2840 ( .A0(n4108), .A1(n8159), .B0(n6878), .B1(n4101), .Y(n5552) );
  OAI22XL U2841 ( .A0(n4190), .A1(n7263), .B0(n6878), .B1(n4183), .Y(n4656) );
  OAI22XL U2842 ( .A0(n4040), .A1(n7520), .B0(n6879), .B1(n5), .Y(n4913) );
  OAI22XL U2843 ( .A0(n4056), .A1(n7648), .B0(n6879), .B1(n6), .Y(n5041) );
  OAI22XL U2844 ( .A0(n4060), .A1(n7776), .B0(n6879), .B1(n4067), .Y(n5169) );
  OAI22XL U2845 ( .A0(n4082), .A1(n7904), .B0(n6879), .B1(n4074), .Y(n5297) );
  OAI22XL U2846 ( .A0(n4094), .A1(n8032), .B0(n6879), .B1(n4087), .Y(n5425) );
  OAI22XL U2847 ( .A0(n4108), .A1(n8160), .B0(n6879), .B1(n4101), .Y(n5553) );
  OAI22XL U2848 ( .A0(n4185), .A1(n7264), .B0(n6879), .B1(n4179), .Y(n4657) );
  OAI22XL U2849 ( .A0(n4043), .A1(n7608), .B0(n6806), .B1(n4038), .Y(n5001) );
  OAI22XL U2850 ( .A0(n4057), .A1(n7736), .B0(n6806), .B1(n4051), .Y(n5129) );
  OAI22XL U2851 ( .A0(n4061), .A1(n7864), .B0(n6806), .B1(n4069), .Y(n5257) );
  OAI22XL U2852 ( .A0(n4082), .A1(n7992), .B0(n6806), .B1(n4079), .Y(n5385) );
  OAI22XL U2853 ( .A0(n6716), .A1(n8120), .B0(n6806), .B1(n4086), .Y(n5513) );
  OAI22XL U2854 ( .A0(n6829), .A1(n8248), .B0(n6806), .B1(n4100), .Y(n5641) );
  OAI22XL U2855 ( .A0(n4189), .A1(n7352), .B0(n6806), .B1(n4182), .Y(n4745) );
  OAI22XL U2856 ( .A0(n4045), .A1(n7609), .B0(n6807), .B1(n4038), .Y(n5002) );
  OAI22XL U2857 ( .A0(n4057), .A1(n7737), .B0(n6807), .B1(n4051), .Y(n5130) );
  OAI22XL U2858 ( .A0(n4060), .A1(n7865), .B0(n6807), .B1(n4069), .Y(n5258) );
  OAI22XL U2859 ( .A0(n4084), .A1(n7993), .B0(n6807), .B1(n4076), .Y(n5386) );
  OAI22XL U2860 ( .A0(n6716), .A1(n8121), .B0(n6807), .B1(n4092), .Y(n5514) );
  OAI22XL U2861 ( .A0(n6829), .A1(n8249), .B0(n6807), .B1(n4106), .Y(n5642) );
  OAI22XL U2862 ( .A0(n4189), .A1(n7353), .B0(n6807), .B1(n4182), .Y(n4746) );
  OAI22XL U2863 ( .A0(n4039), .A1(n7610), .B0(n6808), .B1(n4038), .Y(n5003) );
  OAI22XL U2864 ( .A0(n4057), .A1(n7738), .B0(n6808), .B1(n4051), .Y(n5131) );
  OAI22XL U2865 ( .A0(n4060), .A1(n7866), .B0(n6808), .B1(n4069), .Y(n5259) );
  OAI22XL U2866 ( .A0(n4085), .A1(n7994), .B0(n6808), .B1(n4078), .Y(n5387) );
  OAI22XL U2867 ( .A0(n4099), .A1(n8122), .B0(n6808), .B1(n4086), .Y(n5515) );
  OAI22XL U2868 ( .A0(n4113), .A1(n8250), .B0(n6808), .B1(n4100), .Y(n5643) );
  OAI22XL U2869 ( .A0(n4189), .A1(n7354), .B0(n6808), .B1(n4182), .Y(n4747) );
  OAI22XL U2870 ( .A0(n4041), .A1(n7611), .B0(n6809), .B1(n4034), .Y(n5004) );
  OAI22XL U2871 ( .A0(n4057), .A1(n7739), .B0(n6809), .B1(n4047), .Y(n5132) );
  OAI22XL U2872 ( .A0(n4061), .A1(n7867), .B0(n6809), .B1(n4068), .Y(n5260) );
  OAI22XL U2873 ( .A0(n4081), .A1(n7995), .B0(n6809), .B1(n4075), .Y(n5388) );
  OAI22XL U2874 ( .A0(n4096), .A1(n8123), .B0(n6809), .B1(n4092), .Y(n5516) );
  OAI22XL U2875 ( .A0(n4110), .A1(n8251), .B0(n6809), .B1(n4106), .Y(n5644) );
  OAI22XL U2876 ( .A0(n4189), .A1(n7355), .B0(n6809), .B1(n4182), .Y(n4748) );
  OAI22XL U2877 ( .A0(n4039), .A1(n7612), .B0(n6810), .B1(n4033), .Y(n5005) );
  OAI22XL U2878 ( .A0(n4059), .A1(n7740), .B0(n6810), .B1(n4048), .Y(n5133) );
  OAI22XL U2879 ( .A0(n4062), .A1(n7868), .B0(n6810), .B1(n4068), .Y(n5261) );
  OAI22XL U2880 ( .A0(n4085), .A1(n7996), .B0(n6810), .B1(n4079), .Y(n5389) );
  OAI22XL U2881 ( .A0(n4097), .A1(n8124), .B0(n6810), .B1(n4092), .Y(n5517) );
  OAI22XL U2882 ( .A0(n4111), .A1(n8252), .B0(n6810), .B1(n4106), .Y(n5645) );
  OAI22XL U2883 ( .A0(n4189), .A1(n7356), .B0(n6810), .B1(n4182), .Y(n4749) );
  OAI22XL U2884 ( .A0(n4041), .A1(n7613), .B0(n6811), .B1(n4034), .Y(n5006) );
  OAI22XL U2885 ( .A0(n4053), .A1(n7741), .B0(n6811), .B1(n4047), .Y(n5134) );
  OAI22XL U2886 ( .A0(n4063), .A1(n7869), .B0(n6811), .B1(n4068), .Y(n5262) );
  OAI22XL U2887 ( .A0(n4081), .A1(n7997), .B0(n6811), .B1(n4075), .Y(n5390) );
  OAI22XL U2888 ( .A0(n4095), .A1(n8125), .B0(n6811), .B1(n4092), .Y(n5518) );
  OAI22XL U2889 ( .A0(n4109), .A1(n8253), .B0(n6811), .B1(n4106), .Y(n5646) );
  OAI22XL U2890 ( .A0(n4189), .A1(n7357), .B0(n6811), .B1(n4182), .Y(n4750) );
  OAI22XL U2891 ( .A0(n4040), .A1(n7614), .B0(n6812), .B1(n4038), .Y(n5007) );
  OAI22XL U2892 ( .A0(n4059), .A1(n7742), .B0(n6812), .B1(n4051), .Y(n5135) );
  OAI22XL U2893 ( .A0(n4064), .A1(n7870), .B0(n6812), .B1(n4068), .Y(n5263) );
  OAI22XL U2894 ( .A0(n4085), .A1(n7998), .B0(n6812), .B1(n4076), .Y(n5391) );
  OAI22XL U2895 ( .A0(n4098), .A1(n8126), .B0(n6812), .B1(n4092), .Y(n5519) );
  OAI22XL U2896 ( .A0(n4112), .A1(n8254), .B0(n6812), .B1(n4106), .Y(n5647) );
  OAI22XL U2897 ( .A0(n4189), .A1(n7358), .B0(n6812), .B1(n4182), .Y(n4751) );
  OAI22XL U2898 ( .A0(n4045), .A1(n7615), .B0(n6813), .B1(n5), .Y(n5008) );
  OAI22XL U2899 ( .A0(n4059), .A1(n7743), .B0(n6813), .B1(n4046), .Y(n5136) );
  OAI22XL U2900 ( .A0(n4065), .A1(n7871), .B0(n6813), .B1(n4068), .Y(n5264) );
  OAI22XL U2901 ( .A0(n4081), .A1(n7999), .B0(n6813), .B1(n4075), .Y(n5392) );
  OAI22XL U2902 ( .A0(n4096), .A1(n8127), .B0(n6813), .B1(n4092), .Y(n5520) );
  OAI22XL U2903 ( .A0(n4110), .A1(n8255), .B0(n6813), .B1(n4106), .Y(n5648) );
  OAI22XL U2904 ( .A0(n4189), .A1(n7359), .B0(n6813), .B1(n4182), .Y(n4752) );
  OAI22XL U2905 ( .A0(n4040), .A1(n7616), .B0(n6814), .B1(n4038), .Y(n5009) );
  OAI22XL U2906 ( .A0(n4059), .A1(n7744), .B0(n6814), .B1(n4050), .Y(n5137) );
  OAI22XL U2907 ( .A0(n4065), .A1(n7872), .B0(n6814), .B1(n4068), .Y(n5265) );
  OAI22XL U2908 ( .A0(n4081), .A1(n8000), .B0(n6814), .B1(n4075), .Y(n5393) );
  OAI22XL U2909 ( .A0(n4097), .A1(n8128), .B0(n6814), .B1(n4092), .Y(n5521) );
  OAI22XL U2910 ( .A0(n4111), .A1(n8256), .B0(n6814), .B1(n4106), .Y(n5649) );
  OAI22XL U2911 ( .A0(n4189), .A1(n7360), .B0(n6814), .B1(n4182), .Y(n4753) );
  OAI22XL U2912 ( .A0(n4040), .A1(n7617), .B0(n6815), .B1(n4038), .Y(n5010) );
  OAI22XL U2913 ( .A0(n4059), .A1(n7745), .B0(n6815), .B1(n4049), .Y(n5138) );
  OAI22XL U2914 ( .A0(n4061), .A1(n7873), .B0(n6815), .B1(n4068), .Y(n5266) );
  OAI22XL U2915 ( .A0(n4081), .A1(n8001), .B0(n6815), .B1(n4075), .Y(n5394) );
  OAI22XL U2916 ( .A0(n4095), .A1(n8129), .B0(n6815), .B1(n4092), .Y(n5522) );
  OAI22XL U2917 ( .A0(n4109), .A1(n8257), .B0(n6815), .B1(n4106), .Y(n5650) );
  OAI22XL U2918 ( .A0(n4190), .A1(n7361), .B0(n6815), .B1(n4183), .Y(n4754) );
  OAI22XL U2919 ( .A0(n4040), .A1(n7618), .B0(n6816), .B1(n4038), .Y(n5011) );
  OAI22XL U2920 ( .A0(n4059), .A1(n7746), .B0(n6816), .B1(n4052), .Y(n5139) );
  OAI22XL U2921 ( .A0(n4062), .A1(n7874), .B0(n6816), .B1(n4068), .Y(n5267) );
  OAI22XL U2922 ( .A0(n4082), .A1(n8002), .B0(n6816), .B1(n4075), .Y(n5395) );
  OAI22XL U2923 ( .A0(n4093), .A1(n8130), .B0(n6816), .B1(n4092), .Y(n5523) );
  OAI22XL U2924 ( .A0(n4107), .A1(n8258), .B0(n6816), .B1(n4106), .Y(n5651) );
  OAI22XL U2925 ( .A0(n4190), .A1(n7362), .B0(n6816), .B1(n4183), .Y(n4755) );
  OAI22XL U2926 ( .A0(n4040), .A1(n7619), .B0(n6817), .B1(n4038), .Y(n5012) );
  OAI22XL U2927 ( .A0(n4059), .A1(n7747), .B0(n6817), .B1(n6), .Y(n5140) );
  OAI22XL U2928 ( .A0(n4063), .A1(n7875), .B0(n6817), .B1(n4068), .Y(n5268) );
  OAI22XL U2929 ( .A0(n4084), .A1(n8003), .B0(n6817), .B1(n4075), .Y(n5396) );
  OAI22XL U2930 ( .A0(n4094), .A1(n8131), .B0(n6817), .B1(n4092), .Y(n5524) );
  OAI22XL U2931 ( .A0(n4108), .A1(n8259), .B0(n6817), .B1(n4106), .Y(n5652) );
  OAI22XL U2932 ( .A0(n4190), .A1(n7363), .B0(n6817), .B1(n4183), .Y(n4756) );
  OAI22XL U2933 ( .A0(n4040), .A1(n7620), .B0(n6818), .B1(n4038), .Y(n5013) );
  OAI22XL U2934 ( .A0(n4059), .A1(n7748), .B0(n6818), .B1(n4052), .Y(n5141) );
  OAI22XL U2935 ( .A0(n4064), .A1(n7876), .B0(n6818), .B1(n4068), .Y(n5269) );
  OAI22XL U2936 ( .A0(n4083), .A1(n8004), .B0(n6818), .B1(n4078), .Y(n5397) );
  OAI22XL U2937 ( .A0(n4099), .A1(n8132), .B0(n6818), .B1(n4092), .Y(n5525) );
  OAI22XL U2938 ( .A0(n4113), .A1(n8260), .B0(n6818), .B1(n4106), .Y(n5653) );
  OAI22XL U2939 ( .A0(n4190), .A1(n7364), .B0(n6818), .B1(n4183), .Y(n4757) );
  OAI22XL U2940 ( .A0(n8271), .A1(n6842), .B0(n4352), .B1(n6841), .Y(n4424) );
  AOI2BB1XL U2941 ( .A0N(n7046), .A1N(n4354), .B0(n8289), .Y(n6841) );
  CLKINVX1 U2942 ( .A(n6840), .Y(n4354) );
  OAI22XL U2943 ( .A0(n6720), .A1(n4029), .B0(n6709), .B1(n7394), .Y(n4787) );
  OAI22XL U2944 ( .A0(n6720), .A1(n4067), .B0(n4066), .B1(n7778), .Y(n5171) );
  OAI22XL U2945 ( .A0(n6721), .A1(n4030), .B0(n6709), .B1(n7395), .Y(n4788) );
  OAI22XL U2946 ( .A0(n6721), .A1(n8), .B0(n4066), .B1(n7779), .Y(n5172) );
  OAI22XL U2947 ( .A0(n6722), .A1(n4031), .B0(n6709), .B1(n7396), .Y(n4789) );
  OAI22XL U2948 ( .A0(n6722), .A1(n4072), .B0(n4066), .B1(n7780), .Y(n5173) );
  OAI22XL U2949 ( .A0(n6723), .A1(n4031), .B0(n6709), .B1(n7397), .Y(n4790) );
  OAI22XL U2950 ( .A0(n6723), .A1(n4068), .B0(n4066), .B1(n7781), .Y(n5174) );
  OAI22XL U2951 ( .A0(n6724), .A1(n4025), .B0(n4020), .B1(n7398), .Y(n4791) );
  OAI22XL U2952 ( .A0(n6724), .A1(n4067), .B0(n4066), .B1(n7782), .Y(n5175) );
  OAI22XL U2953 ( .A0(n6725), .A1(n4025), .B0(n4020), .B1(n7399), .Y(n4792) );
  OAI22XL U2954 ( .A0(n6725), .A1(n4070), .B0(n4066), .B1(n7783), .Y(n5176) );
  OAI22XL U2955 ( .A0(n6726), .A1(n4025), .B0(n4020), .B1(n7400), .Y(n4793) );
  OAI22XL U2956 ( .A0(n6726), .A1(n4072), .B0(n4066), .B1(n7784), .Y(n5177) );
  OAI22XL U2957 ( .A0(n6727), .A1(n4025), .B0(n4020), .B1(n7401), .Y(n4794) );
  OAI22XL U2958 ( .A0(n6727), .A1(n4068), .B0(n4066), .B1(n7785), .Y(n5178) );
  OAI22XL U2959 ( .A0(n6728), .A1(n4025), .B0(n4020), .B1(n7402), .Y(n4795) );
  OAI22XL U2960 ( .A0(n6728), .A1(n4071), .B0(n4066), .B1(n7786), .Y(n5179) );
  OAI22XL U2961 ( .A0(n6729), .A1(n4025), .B0(n4021), .B1(n7403), .Y(n4796) );
  OAI22XL U2962 ( .A0(n6729), .A1(n4072), .B0(n4066), .B1(n7787), .Y(n5180) );
  OAI22XL U2963 ( .A0(n6730), .A1(n4025), .B0(n4021), .B1(n7404), .Y(n4797) );
  OAI22XL U2964 ( .A0(n6730), .A1(n4067), .B0(n4066), .B1(n7788), .Y(n5181) );
  OAI22XL U2965 ( .A0(n6731), .A1(n4025), .B0(n4021), .B1(n7405), .Y(n4798) );
  OAI22XL U2966 ( .A0(n6731), .A1(n4068), .B0(n4066), .B1(n7789), .Y(n5182) );
  OAI22XL U2967 ( .A0(n6732), .A1(n4025), .B0(n4021), .B1(n7406), .Y(n4799) );
  OAI22XL U2968 ( .A0(n6732), .A1(n4067), .B0(n6714), .B1(n7790), .Y(n5183) );
  OAI22XL U2969 ( .A0(n6733), .A1(n4025), .B0(n4021), .B1(n7407), .Y(n4800) );
  OAI22XL U2970 ( .A0(n6733), .A1(n4072), .B0(n6714), .B1(n7791), .Y(n5184) );
  OAI22XL U2971 ( .A0(n6734), .A1(n4025), .B0(n4021), .B1(n7408), .Y(n4801) );
  OAI22XL U2972 ( .A0(n6734), .A1(n4068), .B0(n6714), .B1(n7792), .Y(n5185) );
  OAI22XL U2973 ( .A0(n6735), .A1(n4025), .B0(n4021), .B1(n7409), .Y(n4802) );
  OAI22XL U2974 ( .A0(n6735), .A1(n4068), .B0(n6714), .B1(n7793), .Y(n5186) );
  OAI22XL U2975 ( .A0(n6790), .A1(n4030), .B0(n4021), .B1(n7464), .Y(n4857) );
  OAI22XL U2976 ( .A0(n6790), .A1(n4074), .B0(n1334), .B1(n7976), .Y(n5369) );
  OAI22XL U2977 ( .A0(n6791), .A1(n4030), .B0(n4022), .B1(n7465), .Y(n4858) );
  OAI22XL U2978 ( .A0(n6791), .A1(n4074), .B0(n1335), .B1(n7977), .Y(n5370) );
  OAI22XL U2979 ( .A0(n6792), .A1(n4030), .B0(n4023), .B1(n7466), .Y(n4859) );
  OAI22XL U2980 ( .A0(n6792), .A1(n4074), .B0(n1334), .B1(n7978), .Y(n5371) );
  OAI22XL U2981 ( .A0(n6793), .A1(n4030), .B0(n4021), .B1(n7467), .Y(n4860) );
  OAI22XL U2982 ( .A0(n6793), .A1(n4074), .B0(n1335), .B1(n7979), .Y(n5372) );
  OAI22XL U2983 ( .A0(n6794), .A1(n4030), .B0(n4022), .B1(n7468), .Y(n4861) );
  OAI22XL U2984 ( .A0(n6794), .A1(n4080), .B0(n1334), .B1(n7980), .Y(n5373) );
  OAI22XL U2985 ( .A0(n6795), .A1(n4030), .B0(n4023), .B1(n7469), .Y(n4862) );
  OAI22XL U2986 ( .A0(n6795), .A1(n4074), .B0(n1335), .B1(n7981), .Y(n5374) );
  OAI22XL U2987 ( .A0(n6796), .A1(n4030), .B0(n4021), .B1(n7470), .Y(n4863) );
  OAI22XL U2988 ( .A0(n6796), .A1(n4074), .B0(n1334), .B1(n7982), .Y(n5375) );
  OAI22XL U2989 ( .A0(n6862), .A1(n4031), .B0(n4020), .B1(n7375), .Y(n4768) );
  OAI22XL U2990 ( .A0(n6862), .A1(n4080), .B0(n1334), .B1(n7887), .Y(n5280) );
  OAI22XL U2991 ( .A0(n6863), .A1(n4031), .B0(n4020), .B1(n7376), .Y(n4769) );
  OAI22XL U2992 ( .A0(n6863), .A1(n4080), .B0(n1335), .B1(n7888), .Y(n5281) );
  OAI22XL U2993 ( .A0(n6864), .A1(n4029), .B0(n4020), .B1(n7377), .Y(n4770) );
  OAI22XL U2994 ( .A0(n6864), .A1(n4079), .B0(n1334), .B1(n7889), .Y(n5282) );
  OAI22XL U2995 ( .A0(n6865), .A1(n4028), .B0(n4020), .B1(n7378), .Y(n4771) );
  OAI22XL U2996 ( .A0(n6865), .A1(n4079), .B0(n1335), .B1(n7890), .Y(n5283) );
  OAI22XL U2997 ( .A0(n6866), .A1(n4026), .B0(n4020), .B1(n7379), .Y(n4772) );
  OAI22XL U2998 ( .A0(n6866), .A1(n4076), .B0(n1334), .B1(n7891), .Y(n5284) );
  OAI22XL U2999 ( .A0(n6867), .A1(n4027), .B0(n4020), .B1(n7380), .Y(n4773) );
  OAI22XL U3000 ( .A0(n6867), .A1(n4077), .B0(n1335), .B1(n7892), .Y(n5285) );
  OAI22XL U3001 ( .A0(n6797), .A1(n4028), .B0(n4022), .B1(n7471), .Y(n4864) );
  OAI22XL U3002 ( .A0(n6797), .A1(n4074), .B0(n1335), .B1(n7983), .Y(n5376) );
  OAI22XL U3003 ( .A0(n6798), .A1(n4026), .B0(n4023), .B1(n7472), .Y(n4865) );
  OAI22XL U3004 ( .A0(n6798), .A1(n4075), .B0(n1334), .B1(n7984), .Y(n5377) );
  OAI22XL U3005 ( .A0(n6799), .A1(n4027), .B0(n4021), .B1(n7473), .Y(n4866) );
  OAI22XL U3006 ( .A0(n6799), .A1(n4074), .B0(n1335), .B1(n7985), .Y(n5378) );
  OAI22XL U3007 ( .A0(n6800), .A1(n4025), .B0(n4022), .B1(n7474), .Y(n4867) );
  OAI22XL U3008 ( .A0(n6800), .A1(n4074), .B0(n1334), .B1(n7986), .Y(n5379) );
  OAI22XL U3009 ( .A0(n6801), .A1(n4028), .B0(n4023), .B1(n7475), .Y(n4868) );
  OAI22XL U3010 ( .A0(n6801), .A1(n4074), .B0(n1335), .B1(n7987), .Y(n5380) );
  OAI22XL U3011 ( .A0(n6802), .A1(n4025), .B0(n4021), .B1(n7476), .Y(n4869) );
  OAI22XL U3012 ( .A0(n6802), .A1(n4079), .B0(n1334), .B1(n7988), .Y(n5381) );
  OAI22XL U3013 ( .A0(n6803), .A1(n4030), .B0(n4022), .B1(n7477), .Y(n4870) );
  OAI22XL U3014 ( .A0(n6803), .A1(n4079), .B0(n1335), .B1(n7989), .Y(n5382) );
  OAI22XL U3015 ( .A0(n6804), .A1(n4030), .B0(n4023), .B1(n7478), .Y(n4871) );
  OAI22XL U3016 ( .A0(n6804), .A1(n4078), .B0(n1334), .B1(n7990), .Y(n5383) );
  OAI22XL U3017 ( .A0(n6805), .A1(n4026), .B0(n4021), .B1(n7479), .Y(n4872) );
  OAI22XL U3018 ( .A0(n6805), .A1(n4074), .B0(n1335), .B1(n7991), .Y(n5384) );
  OAI22XL U3019 ( .A0(n6819), .A1(n4029), .B0(n4019), .B1(n7493), .Y(n4886) );
  OAI22XL U3020 ( .A0(n6819), .A1(n4067), .B0(n6714), .B1(n7877), .Y(n5270) );
  OAI22XL U3021 ( .A0(n6820), .A1(n4026), .B0(n4019), .B1(n7494), .Y(n4887) );
  OAI22XL U3022 ( .A0(n6820), .A1(n4067), .B0(n6714), .B1(n7878), .Y(n5271) );
  OAI22XL U3023 ( .A0(n6821), .A1(n7), .B0(n6709), .B1(n7495), .Y(n4888) );
  OAI22XL U3024 ( .A0(n6821), .A1(n4067), .B0(n6714), .B1(n7879), .Y(n5272) );
  OAI22XL U3025 ( .A0(n6822), .A1(n7), .B0(n6709), .B1(n7496), .Y(n4889) );
  OAI22XL U3026 ( .A0(n6822), .A1(n4067), .B0(n6714), .B1(n7880), .Y(n5273) );
  OAI22XL U3027 ( .A0(n6823), .A1(n4028), .B0(n4022), .B1(n7497), .Y(n4890) );
  OAI22XL U3028 ( .A0(n6823), .A1(n4067), .B0(n6714), .B1(n7881), .Y(n5274) );
  OAI22XL U3029 ( .A0(n6824), .A1(n4029), .B0(n4023), .B1(n7498), .Y(n4891) );
  OAI22XL U3030 ( .A0(n6824), .A1(n4067), .B0(n6714), .B1(n7882), .Y(n5275) );
  OAI22XL U3031 ( .A0(n6825), .A1(n4029), .B0(n4021), .B1(n7499), .Y(n4892) );
  OAI22XL U3032 ( .A0(n6825), .A1(n4067), .B0(n6714), .B1(n7883), .Y(n5276) );
  OAI22XL U3033 ( .A0(n6826), .A1(n4031), .B0(n4022), .B1(n7500), .Y(n4893) );
  OAI22XL U3034 ( .A0(n6826), .A1(n4067), .B0(n6714), .B1(n7884), .Y(n5277) );
  OAI22XL U3035 ( .A0(n6827), .A1(n4031), .B0(n4022), .B1(n7501), .Y(n4894) );
  OAI22XL U3036 ( .A0(n6827), .A1(n4067), .B0(n4066), .B1(n7885), .Y(n5278) );
  OAI22XL U3037 ( .A0(n6828), .A1(n4028), .B0(n4023), .B1(n7502), .Y(n4895) );
  OAI22XL U3038 ( .A0(n6828), .A1(n4068), .B0(n4066), .B1(n7886), .Y(n5279) );
  OAI22XL U3039 ( .A0(n6719), .A1(n4026), .B0(n4019), .B1(n7393), .Y(n4786) );
  OAI22XL U3040 ( .A0(n6736), .A1(n4025), .B0(n4021), .B1(n7410), .Y(n4803) );
  OAI22XL U3041 ( .A0(n6737), .A1(n4026), .B0(n4021), .B1(n7411), .Y(n4804) );
  OAI22XL U3042 ( .A0(n6738), .A1(n4026), .B0(n4021), .B1(n7412), .Y(n4805) );
  OAI22XL U3043 ( .A0(n6739), .A1(n4026), .B0(n4021), .B1(n7413), .Y(n4806) );
  OAI22XL U3044 ( .A0(n6740), .A1(n4026), .B0(n4021), .B1(n7414), .Y(n4807) );
  OAI22XL U3045 ( .A0(n6741), .A1(n4026), .B0(n4022), .B1(n7415), .Y(n4808) );
  OAI22XL U3046 ( .A0(n6742), .A1(n4026), .B0(n4022), .B1(n7416), .Y(n4809) );
  OAI22XL U3047 ( .A0(n6743), .A1(n4026), .B0(n4022), .B1(n7417), .Y(n4810) );
  OAI22XL U3048 ( .A0(n6744), .A1(n4026), .B0(n4022), .B1(n7418), .Y(n4811) );
  OAI22XL U3049 ( .A0(n6745), .A1(n4026), .B0(n4022), .B1(n7419), .Y(n4812) );
  OAI22XL U3050 ( .A0(n6746), .A1(n4026), .B0(n4022), .B1(n7420), .Y(n4813) );
  OAI22XL U3051 ( .A0(n6747), .A1(n4026), .B0(n4022), .B1(n7421), .Y(n4814) );
  OAI22XL U3052 ( .A0(n6748), .A1(n4026), .B0(n4022), .B1(n7422), .Y(n4815) );
  OAI22XL U3053 ( .A0(n6749), .A1(n4027), .B0(n4022), .B1(n7423), .Y(n4816) );
  OAI22XL U3054 ( .A0(n6750), .A1(n4027), .B0(n4022), .B1(n7424), .Y(n4817) );
  OAI22XL U3055 ( .A0(n6751), .A1(n4027), .B0(n4022), .B1(n7425), .Y(n4818) );
  OAI22XL U3056 ( .A0(n6752), .A1(n4027), .B0(n4022), .B1(n7426), .Y(n4819) );
  OAI22XL U3057 ( .A0(n6753), .A1(n4027), .B0(n4023), .B1(n7427), .Y(n4820) );
  OAI22XL U3058 ( .A0(n6754), .A1(n4027), .B0(n4023), .B1(n7428), .Y(n4821) );
  OAI22XL U3059 ( .A0(n6755), .A1(n4027), .B0(n4023), .B1(n7429), .Y(n4822) );
  OAI22XL U3060 ( .A0(n6756), .A1(n4027), .B0(n4023), .B1(n7430), .Y(n4823) );
  OAI22XL U3061 ( .A0(n6757), .A1(n4027), .B0(n4023), .B1(n7431), .Y(n4824) );
  OAI22XL U3062 ( .A0(n6758), .A1(n4027), .B0(n4023), .B1(n7432), .Y(n4825) );
  OAI22XL U3063 ( .A0(n6759), .A1(n4027), .B0(n4023), .B1(n7433), .Y(n4826) );
  OAI22XL U3064 ( .A0(n6760), .A1(n4027), .B0(n4023), .B1(n7434), .Y(n4827) );
  OAI22XL U3065 ( .A0(n6761), .A1(n4028), .B0(n4023), .B1(n7435), .Y(n4828) );
  OAI22XL U3066 ( .A0(n6762), .A1(n4028), .B0(n4023), .B1(n7436), .Y(n4829) );
  OAI22XL U3067 ( .A0(n6763), .A1(n4028), .B0(n4023), .B1(n7437), .Y(n4830) );
  OAI22XL U3068 ( .A0(n6764), .A1(n4028), .B0(n4023), .B1(n7438), .Y(n4831) );
  OAI22XL U3069 ( .A0(n6765), .A1(n4028), .B0(n4021), .B1(n7439), .Y(n4832) );
  OAI22XL U3070 ( .A0(n6766), .A1(n4028), .B0(n4023), .B1(n7440), .Y(n4833) );
  OAI22XL U3071 ( .A0(n6767), .A1(n4028), .B0(n4022), .B1(n7441), .Y(n4834) );
  OAI22XL U3072 ( .A0(n6768), .A1(n4028), .B0(n4024), .B1(n7442), .Y(n4835) );
  OAI22XL U3073 ( .A0(n6769), .A1(n4028), .B0(n4020), .B1(n7443), .Y(n4836) );
  OAI22XL U3074 ( .A0(n6770), .A1(n4028), .B0(n4020), .B1(n7444), .Y(n4837) );
  OAI22XL U3075 ( .A0(n6771), .A1(n4028), .B0(n6710), .B1(n7445), .Y(n4838) );
  OAI22XL U3076 ( .A0(n6772), .A1(n4028), .B0(n6710), .B1(n7446), .Y(n4839) );
  OAI22XL U3077 ( .A0(n6773), .A1(n4029), .B0(n4020), .B1(n7447), .Y(n4840) );
  OAI22XL U3078 ( .A0(n6774), .A1(n4029), .B0(n4020), .B1(n7448), .Y(n4841) );
  OAI22XL U3079 ( .A0(n6775), .A1(n4029), .B0(n4020), .B1(n7449), .Y(n4842) );
  OAI22XL U3080 ( .A0(n6776), .A1(n4029), .B0(n4020), .B1(n7450), .Y(n4843) );
  OAI22XL U3081 ( .A0(n6777), .A1(n4029), .B0(n4024), .B1(n7451), .Y(n4844) );
  OAI22XL U3082 ( .A0(n6778), .A1(n4029), .B0(n4024), .B1(n7452), .Y(n4845) );
  OAI22XL U3083 ( .A0(n6779), .A1(n4029), .B0(n4024), .B1(n7453), .Y(n4846) );
  OAI22XL U3084 ( .A0(n6780), .A1(n4029), .B0(n4024), .B1(n7454), .Y(n4847) );
  OAI22XL U3085 ( .A0(n6781), .A1(n4029), .B0(n4024), .B1(n7455), .Y(n4848) );
  OAI22XL U3086 ( .A0(n6782), .A1(n4029), .B0(n4024), .B1(n7456), .Y(n4849) );
  OAI22XL U3087 ( .A0(n6783), .A1(n4029), .B0(n4024), .B1(n7457), .Y(n4850) );
  OAI22XL U3088 ( .A0(n6784), .A1(n4029), .B0(n4024), .B1(n7458), .Y(n4851) );
  OAI22XL U3089 ( .A0(n6785), .A1(n4030), .B0(n4024), .B1(n7459), .Y(n4852) );
  OAI22XL U3090 ( .A0(n6786), .A1(n4030), .B0(n4024), .B1(n7460), .Y(n4853) );
  OAI22XL U3091 ( .A0(n6787), .A1(n4030), .B0(n4024), .B1(n7461), .Y(n4854) );
  OAI22XL U3092 ( .A0(n6788), .A1(n4030), .B0(n4024), .B1(n7462), .Y(n4855) );
  OAI22XL U3093 ( .A0(n6789), .A1(n4030), .B0(n4023), .B1(n7463), .Y(n4856) );
  OAI22XL U3094 ( .A0(n6868), .A1(n4025), .B0(n4020), .B1(n7381), .Y(n4774) );
  OAI22XL U3095 ( .A0(n6869), .A1(n4027), .B0(n4019), .B1(n7382), .Y(n4775) );
  OAI22XL U3096 ( .A0(n6870), .A1(n4025), .B0(n4019), .B1(n7383), .Y(n4776) );
  OAI22XL U3097 ( .A0(n6871), .A1(n4030), .B0(n4019), .B1(n7384), .Y(n4777) );
  OAI22XL U3098 ( .A0(n6872), .A1(n4031), .B0(n4019), .B1(n7385), .Y(n4778) );
  OAI22XL U3099 ( .A0(n6873), .A1(n4031), .B0(n4019), .B1(n7386), .Y(n4779) );
  OAI22XL U3100 ( .A0(n6874), .A1(n4027), .B0(n4019), .B1(n7387), .Y(n4780) );
  OAI22XL U3101 ( .A0(n6875), .A1(n4025), .B0(n4019), .B1(n7388), .Y(n4781) );
  OAI22XL U3102 ( .A0(n6876), .A1(n4030), .B0(n4019), .B1(n7389), .Y(n4782) );
  OAI22XL U3103 ( .A0(n6877), .A1(n4028), .B0(n4019), .B1(n7390), .Y(n4783) );
  OAI22XL U3104 ( .A0(n6878), .A1(n4026), .B0(n4019), .B1(n7391), .Y(n4784) );
  OAI22XL U3105 ( .A0(n6879), .A1(n4027), .B0(n4019), .B1(n7392), .Y(n4785) );
  OAI22XL U3106 ( .A0(n6806), .A1(n4027), .B0(n4021), .B1(n7480), .Y(n4873) );
  OAI22XL U3107 ( .A0(n6807), .A1(n4030), .B0(n6709), .B1(n7481), .Y(n4874) );
  OAI22XL U3108 ( .A0(n6808), .A1(n4031), .B0(n6709), .B1(n7482), .Y(n4875) );
  OAI22XL U3109 ( .A0(n6809), .A1(n7), .B0(n6709), .B1(n7483), .Y(n4876) );
  OAI22XL U3110 ( .A0(n6810), .A1(n4029), .B0(n4019), .B1(n7484), .Y(n4877) );
  OAI22XL U3111 ( .A0(n6811), .A1(n4031), .B0(n4019), .B1(n7485), .Y(n4878) );
  OAI22XL U3112 ( .A0(n6812), .A1(n4031), .B0(n4019), .B1(n7486), .Y(n4879) );
  OAI22XL U3113 ( .A0(n6813), .A1(n7), .B0(n4019), .B1(n7487), .Y(n4880) );
  OAI22XL U3114 ( .A0(n6814), .A1(n7), .B0(n4019), .B1(n7488), .Y(n4881) );
  OAI22XL U3115 ( .A0(n6815), .A1(n7), .B0(n6709), .B1(n7489), .Y(n4882) );
  OAI22XL U3116 ( .A0(n6816), .A1(n4031), .B0(n6709), .B1(n7490), .Y(n4883) );
  OAI22XL U3117 ( .A0(n6817), .A1(n4031), .B0(n6709), .B1(n7491), .Y(n4884) );
  OAI22XL U3118 ( .A0(n6818), .A1(n4031), .B0(n6709), .B1(n7492), .Y(n4885) );
  CLKBUFX3 U3119 ( .A(n6718), .Y(n1333) );
  AOI211XL U3120 ( .A0(n4421), .A1(n1345), .B0(n4353), .C0(n8289), .Y(n6718)
         );
  CLKINVX1 U3121 ( .A(n6843), .Y(n4353) );
  NAND3X2 U3122 ( .A(n7045), .B(n8272), .C(n6843), .Y(n6844) );
  NOR4X1 U3123 ( .A(n6836), .B(n6835), .C(n6834), .D(n6833), .Y(n6840) );
  OAI22XL U3124 ( .A0(n4135), .A1(n8287), .B0(n4145), .B1(n8288), .Y(n6834) );
  OAI22XL U3125 ( .A0(n4115), .A1(n8285), .B0(n4125), .B1(n8286), .Y(n6833) );
  OAI22XL U3126 ( .A0(n1697), .A1(n8283), .B0(n1355), .B1(n8284), .Y(n6836) );
  OAI22XL U3127 ( .A0(n4175), .A1(n7048), .B0(n4397), .B1(n4177), .Y(n4616) );
  OAI22XL U3128 ( .A0(n1295), .A1(n7049), .B0(n4398), .B1(n6861), .Y(n4617) );
  OAI22XL U3129 ( .A0(n4175), .A1(n7050), .B0(n4399), .B1(n4176), .Y(n4618) );
  OAI22XL U3130 ( .A0(n4175), .A1(n7051), .B0(n4400), .B1(n4177), .Y(n4619) );
  OAI22XL U3131 ( .A0(n4175), .A1(n7052), .B0(n4401), .B1(n4176), .Y(n4620) );
  OAI22XL U3132 ( .A0(n4175), .A1(n7053), .B0(n4402), .B1(n4176), .Y(n4621) );
  OAI22XL U3133 ( .A0(n4175), .A1(n7054), .B0(n4403), .B1(n4176), .Y(n4622) );
  OAI22XL U3134 ( .A0(n4175), .A1(n7055), .B0(n4404), .B1(n4176), .Y(n4623) );
  OAI22XL U3135 ( .A0(n4175), .A1(n7056), .B0(n4405), .B1(n4176), .Y(n4624) );
  OAI22XL U3136 ( .A0(n4175), .A1(n7057), .B0(n4406), .B1(n4176), .Y(n4625) );
  OAI22XL U3137 ( .A0(n1295), .A1(n7058), .B0(n4407), .B1(n4176), .Y(n4626) );
  OAI22XL U3138 ( .A0(n4175), .A1(n7059), .B0(n4408), .B1(n4177), .Y(n4627) );
  OAI22XL U3139 ( .A0(n4175), .A1(n7060), .B0(n4409), .B1(n6861), .Y(n4628) );
  OAI22XL U3140 ( .A0(n4175), .A1(n7061), .B0(n4410), .B1(n4176), .Y(n4629) );
  OAI22XL U3141 ( .A0(n4175), .A1(n7062), .B0(n4411), .B1(n4177), .Y(n4630) );
  OAI22XL U3142 ( .A0(n4175), .A1(n7063), .B0(n4412), .B1(n4177), .Y(n4631) );
  OAI22XL U3143 ( .A0(n4175), .A1(n7064), .B0(n4413), .B1(n4177), .Y(n4632) );
  OAI22XL U3144 ( .A0(n4175), .A1(n7065), .B0(n4414), .B1(n4176), .Y(n4633) );
  OAI22XL U3145 ( .A0(n4175), .A1(n7066), .B0(n4415), .B1(n4177), .Y(n4634) );
  OAI22XL U3146 ( .A0(n4175), .A1(n7067), .B0(n4416), .B1(n4177), .Y(n4635) );
  OAI22XL U3147 ( .A0(n4175), .A1(n7068), .B0(n4417), .B1(n4177), .Y(n4636) );
  OAI22XL U3148 ( .A0(n4175), .A1(n7069), .B0(n4418), .B1(n4177), .Y(n4637) );
  OAI22XL U3149 ( .A0(n4175), .A1(n7070), .B0(n4419), .B1(n4177), .Y(n4638) );
  OAI2BB2XL U3150 ( .B0(n4420), .B1(n4177), .A0N(n4176), .A1N(n1297), .Y(n4639) );
  OAI22XL U3151 ( .A0(n4154), .A1(n7222), .B0(n4396), .B1(n4156), .Y(n4441) );
  OAI22XL U3152 ( .A0(n4154), .A1(n7223), .B0(n4397), .B1(n4155), .Y(n4442) );
  OAI22XL U3153 ( .A0(n4154), .A1(n7224), .B0(n4398), .B1(n6850), .Y(n4443) );
  OAI22XL U3154 ( .A0(n4154), .A1(n7225), .B0(n4399), .B1(n4155), .Y(n4444) );
  OAI22XL U3155 ( .A0(n4154), .A1(n7226), .B0(n4400), .B1(n4156), .Y(n4445) );
  OAI22XL U3156 ( .A0(n4154), .A1(n7227), .B0(n4401), .B1(n4155), .Y(n4446) );
  OAI22XL U3157 ( .A0(n4154), .A1(n7228), .B0(n4402), .B1(n4155), .Y(n4447) );
  OAI22XL U3158 ( .A0(n4154), .A1(n7229), .B0(n4403), .B1(n4155), .Y(n4448) );
  OAI22XL U3159 ( .A0(n4154), .A1(n7230), .B0(n4404), .B1(n4155), .Y(n4449) );
  OAI22XL U3160 ( .A0(n4154), .A1(n7231), .B0(n4405), .B1(n4155), .Y(n4450) );
  OAI22XL U3161 ( .A0(n4154), .A1(n7232), .B0(n4406), .B1(n4155), .Y(n4451) );
  OAI22XL U3162 ( .A0(n4154), .A1(n7233), .B0(n4407), .B1(n4155), .Y(n4452) );
  OAI22XL U3163 ( .A0(n4154), .A1(n7234), .B0(n4408), .B1(n4156), .Y(n4453) );
  OAI22XL U3164 ( .A0(n1289), .A1(n7235), .B0(n4409), .B1(n6850), .Y(n4454) );
  OAI22XL U3165 ( .A0(n1289), .A1(n7236), .B0(n4410), .B1(n4155), .Y(n4455) );
  OAI22XL U3166 ( .A0(n4154), .A1(n7237), .B0(n4411), .B1(n4156), .Y(n4456) );
  OAI22XL U3167 ( .A0(n4154), .A1(n7238), .B0(n4412), .B1(n4156), .Y(n4457) );
  OAI22XL U3168 ( .A0(n4154), .A1(n7239), .B0(n4413), .B1(n4156), .Y(n4458) );
  OAI22XL U3169 ( .A0(n1289), .A1(n7240), .B0(n4414), .B1(n4155), .Y(n4459) );
  OAI22XL U3170 ( .A0(n4154), .A1(n7241), .B0(n4415), .B1(n4156), .Y(n4460) );
  OAI22XL U3171 ( .A0(n4154), .A1(n7242), .B0(n4416), .B1(n4156), .Y(n4461) );
  OAI22XL U3172 ( .A0(n4154), .A1(n7243), .B0(n4417), .B1(n4156), .Y(n4462) );
  OAI22XL U3173 ( .A0(n4154), .A1(n7244), .B0(n4418), .B1(n4156), .Y(n4463) );
  OAI22XL U3174 ( .A0(n4154), .A1(n7245), .B0(n4419), .B1(n4156), .Y(n4464) );
  OAI2BB2XL U3175 ( .B0(n4420), .B1(n4156), .A0N(n4155), .A1N(n1298), .Y(n4465) );
  OAI22XL U3176 ( .A0(n4157), .A1(n7197), .B0(n4396), .B1(n4159), .Y(n4466) );
  OAI22XL U3177 ( .A0(n4157), .A1(n7198), .B0(n4397), .B1(n4158), .Y(n4467) );
  OAI22XL U3178 ( .A0(n4157), .A1(n7199), .B0(n4398), .B1(n6851), .Y(n4468) );
  OAI22XL U3179 ( .A0(n4157), .A1(n7200), .B0(n4399), .B1(n4158), .Y(n4469) );
  OAI22XL U3180 ( .A0(n4157), .A1(n7201), .B0(n4400), .B1(n4159), .Y(n4470) );
  OAI22XL U3181 ( .A0(n4157), .A1(n7202), .B0(n4401), .B1(n4158), .Y(n4471) );
  OAI22XL U3182 ( .A0(n4157), .A1(n7203), .B0(n4402), .B1(n4158), .Y(n4472) );
  OAI22XL U3183 ( .A0(n4157), .A1(n7204), .B0(n4403), .B1(n4158), .Y(n4473) );
  OAI22XL U3184 ( .A0(n4157), .A1(n7205), .B0(n4404), .B1(n4158), .Y(n4474) );
  OAI22XL U3185 ( .A0(n4157), .A1(n7206), .B0(n4405), .B1(n4158), .Y(n4475) );
  OAI22XL U3186 ( .A0(n4157), .A1(n7207), .B0(n4406), .B1(n4158), .Y(n4476) );
  OAI22XL U3187 ( .A0(n4157), .A1(n7208), .B0(n4407), .B1(n4158), .Y(n4477) );
  OAI22XL U3188 ( .A0(n4157), .A1(n7209), .B0(n4408), .B1(n4159), .Y(n4478) );
  OAI22XL U3189 ( .A0(n1290), .A1(n7210), .B0(n4409), .B1(n6851), .Y(n4479) );
  OAI22XL U3190 ( .A0(n1290), .A1(n7211), .B0(n4410), .B1(n4158), .Y(n4480) );
  OAI22XL U3191 ( .A0(n4157), .A1(n7212), .B0(n4411), .B1(n4159), .Y(n4481) );
  OAI22XL U3192 ( .A0(n4157), .A1(n7213), .B0(n4412), .B1(n4159), .Y(n4482) );
  OAI22XL U3193 ( .A0(n4157), .A1(n7214), .B0(n4413), .B1(n4159), .Y(n4483) );
  OAI22XL U3194 ( .A0(n1290), .A1(n7215), .B0(n4414), .B1(n4158), .Y(n4484) );
  OAI22XL U3195 ( .A0(n4157), .A1(n7216), .B0(n4415), .B1(n4159), .Y(n4485) );
  OAI22XL U3196 ( .A0(n4157), .A1(n7217), .B0(n4416), .B1(n4159), .Y(n4486) );
  OAI22XL U3197 ( .A0(n4157), .A1(n7218), .B0(n4417), .B1(n4159), .Y(n4487) );
  OAI22XL U3198 ( .A0(n4157), .A1(n7219), .B0(n4418), .B1(n4159), .Y(n4488) );
  OAI22XL U3199 ( .A0(n4157), .A1(n7220), .B0(n4419), .B1(n4159), .Y(n4489) );
  OAI2BB2XL U3200 ( .B0(n4420), .B1(n4159), .A0N(n4158), .A1N(n1299), .Y(n4490) );
  OAI22XL U3201 ( .A0(n4160), .A1(n7172), .B0(n4396), .B1(n4162), .Y(n4491) );
  OAI22XL U3202 ( .A0(n4160), .A1(n7173), .B0(n4397), .B1(n4161), .Y(n4492) );
  OAI22XL U3203 ( .A0(n4160), .A1(n7174), .B0(n4398), .B1(n6852), .Y(n4493) );
  OAI22XL U3204 ( .A0(n4160), .A1(n7175), .B0(n4399), .B1(n4161), .Y(n4494) );
  OAI22XL U3205 ( .A0(n4160), .A1(n7176), .B0(n4400), .B1(n4162), .Y(n4495) );
  OAI22XL U3206 ( .A0(n4160), .A1(n7177), .B0(n4401), .B1(n4161), .Y(n4496) );
  OAI22XL U3207 ( .A0(n4160), .A1(n7178), .B0(n4402), .B1(n4161), .Y(n4497) );
  OAI22XL U3208 ( .A0(n4160), .A1(n7179), .B0(n4403), .B1(n4161), .Y(n4498) );
  OAI22XL U3209 ( .A0(n4160), .A1(n7180), .B0(n4404), .B1(n4161), .Y(n4499) );
  OAI22XL U3210 ( .A0(n4160), .A1(n7181), .B0(n4405), .B1(n4161), .Y(n4500) );
  OAI22XL U3211 ( .A0(n4160), .A1(n7182), .B0(n4406), .B1(n4161), .Y(n4501) );
  OAI22XL U3212 ( .A0(n4160), .A1(n7183), .B0(n4407), .B1(n4161), .Y(n4502) );
  OAI22XL U3213 ( .A0(n4160), .A1(n7184), .B0(n4408), .B1(n4162), .Y(n4503) );
  OAI22XL U3214 ( .A0(n1291), .A1(n7185), .B0(n4409), .B1(n6852), .Y(n4504) );
  OAI22XL U3215 ( .A0(n1291), .A1(n7186), .B0(n4410), .B1(n4161), .Y(n4505) );
  OAI22XL U3216 ( .A0(n4160), .A1(n7187), .B0(n4411), .B1(n4162), .Y(n4506) );
  OAI22XL U3217 ( .A0(n4160), .A1(n7188), .B0(n4412), .B1(n4162), .Y(n4507) );
  OAI22XL U3218 ( .A0(n4160), .A1(n7189), .B0(n4413), .B1(n4162), .Y(n4508) );
  OAI22XL U3219 ( .A0(n1291), .A1(n7190), .B0(n4414), .B1(n4161), .Y(n4509) );
  OAI22XL U3220 ( .A0(n4160), .A1(n7191), .B0(n4415), .B1(n4162), .Y(n4510) );
  OAI22XL U3221 ( .A0(n4160), .A1(n7192), .B0(n4416), .B1(n4162), .Y(n4511) );
  OAI22XL U3222 ( .A0(n4160), .A1(n7193), .B0(n4417), .B1(n4162), .Y(n4512) );
  OAI22XL U3223 ( .A0(n4160), .A1(n7194), .B0(n4418), .B1(n4162), .Y(n4513) );
  OAI22XL U3224 ( .A0(n4160), .A1(n7195), .B0(n4419), .B1(n4162), .Y(n4514) );
  OAI22XL U3225 ( .A0(n4163), .A1(n7147), .B0(n4396), .B1(n4164), .Y(n4516) );
  OAI22XL U3226 ( .A0(n4163), .A1(n7148), .B0(n4397), .B1(n4164), .Y(n4517) );
  OAI22XL U3227 ( .A0(n4163), .A1(n7149), .B0(n4398), .B1(n4164), .Y(n4518) );
  OAI22XL U3228 ( .A0(n4163), .A1(n7150), .B0(n4399), .B1(n4165), .Y(n4519) );
  OAI22XL U3229 ( .A0(n4163), .A1(n7151), .B0(n4400), .B1(n4165), .Y(n4520) );
  OAI22XL U3230 ( .A0(n4163), .A1(n7152), .B0(n4401), .B1(n4165), .Y(n4521) );
  OAI22XL U3231 ( .A0(n4163), .A1(n7153), .B0(n4402), .B1(n4164), .Y(n4522) );
  OAI22XL U3232 ( .A0(n4163), .A1(n7154), .B0(n4403), .B1(n6853), .Y(n4523) );
  OAI22XL U3233 ( .A0(n4163), .A1(n7155), .B0(n4404), .B1(n6853), .Y(n4524) );
  OAI22XL U3234 ( .A0(n4163), .A1(n7156), .B0(n4405), .B1(n4165), .Y(n4525) );
  OAI22XL U3235 ( .A0(n4163), .A1(n7157), .B0(n4406), .B1(n4164), .Y(n4526) );
  OAI22XL U3236 ( .A0(n4163), .A1(n7158), .B0(n4407), .B1(n4165), .Y(n4527) );
  OAI22XL U3237 ( .A0(n4163), .A1(n7159), .B0(n4408), .B1(n4165), .Y(n4528) );
  OAI22XL U3238 ( .A0(n4163), .A1(n7160), .B0(n4409), .B1(n4165), .Y(n4529) );
  OAI22XL U3239 ( .A0(n4163), .A1(n7161), .B0(n4410), .B1(n4165), .Y(n4530) );
  OAI22XL U3240 ( .A0(n4163), .A1(n7162), .B0(n4411), .B1(n4165), .Y(n4531) );
  OAI22XL U3241 ( .A0(n4163), .A1(n7163), .B0(n4412), .B1(n4165), .Y(n4532) );
  OAI22XL U3242 ( .A0(n4163), .A1(n7164), .B0(n4413), .B1(n4164), .Y(n4533) );
  OAI22XL U3243 ( .A0(n4163), .A1(n7165), .B0(n4414), .B1(n4164), .Y(n4534) );
  OAI22XL U3244 ( .A0(n4163), .A1(n7166), .B0(n4415), .B1(n4165), .Y(n4535) );
  OAI22XL U3245 ( .A0(n4163), .A1(n7167), .B0(n4416), .B1(n4164), .Y(n4536) );
  OAI22XL U3246 ( .A0(n1292), .A1(n7168), .B0(n4417), .B1(n4164), .Y(n4537) );
  OAI22XL U3247 ( .A0(n1292), .A1(n7169), .B0(n4418), .B1(n4164), .Y(n4538) );
  OAI22XL U3248 ( .A0(n1292), .A1(n7170), .B0(n4419), .B1(n4164), .Y(n4539) );
  OAI22XL U3249 ( .A0(n4166), .A1(n7122), .B0(n4396), .B1(n4168), .Y(n4541) );
  OAI22XL U3250 ( .A0(n4166), .A1(n7123), .B0(n4397), .B1(n4167), .Y(n4542) );
  OAI22XL U3251 ( .A0(n4166), .A1(n7124), .B0(n4398), .B1(n6855), .Y(n4543) );
  OAI22XL U3252 ( .A0(n4166), .A1(n7125), .B0(n4399), .B1(n4167), .Y(n4544) );
  OAI22XL U3253 ( .A0(n4166), .A1(n7126), .B0(n4400), .B1(n4168), .Y(n4545) );
  OAI22XL U3254 ( .A0(n4166), .A1(n7127), .B0(n4401), .B1(n4167), .Y(n4546) );
  OAI22XL U3255 ( .A0(n4166), .A1(n7128), .B0(n4402), .B1(n4167), .Y(n4547) );
  OAI22XL U3256 ( .A0(n4166), .A1(n7129), .B0(n4403), .B1(n4167), .Y(n4548) );
  OAI22XL U3257 ( .A0(n4166), .A1(n7130), .B0(n4404), .B1(n4167), .Y(n4549) );
  OAI22XL U3258 ( .A0(n4166), .A1(n7131), .B0(n4405), .B1(n4167), .Y(n4550) );
  OAI22XL U3259 ( .A0(n4166), .A1(n7132), .B0(n4406), .B1(n4167), .Y(n4551) );
  OAI22XL U3260 ( .A0(n4166), .A1(n7133), .B0(n4407), .B1(n4167), .Y(n4552) );
  OAI22XL U3261 ( .A0(n4166), .A1(n7134), .B0(n4408), .B1(n4168), .Y(n4553) );
  OAI22XL U3262 ( .A0(n1293), .A1(n7135), .B0(n4409), .B1(n6855), .Y(n4554) );
  OAI22XL U3263 ( .A0(n1293), .A1(n7136), .B0(n4410), .B1(n4167), .Y(n4555) );
  OAI22XL U3264 ( .A0(n4166), .A1(n7137), .B0(n4411), .B1(n4168), .Y(n4556) );
  OAI22XL U3265 ( .A0(n4166), .A1(n7138), .B0(n4412), .B1(n4168), .Y(n4557) );
  OAI22XL U3266 ( .A0(n4166), .A1(n7139), .B0(n4413), .B1(n4168), .Y(n4558) );
  OAI22XL U3267 ( .A0(n1293), .A1(n7140), .B0(n4414), .B1(n4167), .Y(n4559) );
  OAI22XL U3268 ( .A0(n4166), .A1(n7141), .B0(n4415), .B1(n4168), .Y(n4560) );
  OAI22XL U3269 ( .A0(n4166), .A1(n7142), .B0(n4416), .B1(n4168), .Y(n4561) );
  OAI22XL U3270 ( .A0(n4166), .A1(n7143), .B0(n4417), .B1(n4168), .Y(n4562) );
  OAI22XL U3271 ( .A0(n4166), .A1(n7144), .B0(n4418), .B1(n4168), .Y(n4563) );
  OAI22XL U3272 ( .A0(n4166), .A1(n7145), .B0(n4419), .B1(n4168), .Y(n4564) );
  OAI2BB2XL U3273 ( .B0(n4420), .B1(n4168), .A0N(n4167), .A1N(n1300), .Y(n4565) );
  OAI22XL U3274 ( .A0(n4169), .A1(n7097), .B0(n4396), .B1(n4171), .Y(n4566) );
  OAI22XL U3275 ( .A0(n4169), .A1(n7098), .B0(n4397), .B1(n4170), .Y(n4567) );
  OAI22XL U3276 ( .A0(n4169), .A1(n7099), .B0(n4398), .B1(n6857), .Y(n4568) );
  OAI22XL U3277 ( .A0(n4169), .A1(n7100), .B0(n4399), .B1(n4170), .Y(n4569) );
  OAI22XL U3278 ( .A0(n4169), .A1(n7101), .B0(n4400), .B1(n4171), .Y(n4570) );
  OAI22XL U3279 ( .A0(n4169), .A1(n7102), .B0(n4401), .B1(n4170), .Y(n4571) );
  OAI22XL U3280 ( .A0(n4169), .A1(n7103), .B0(n4402), .B1(n4170), .Y(n4572) );
  OAI22XL U3281 ( .A0(n4169), .A1(n7104), .B0(n4403), .B1(n4170), .Y(n4573) );
  OAI22XL U3282 ( .A0(n4169), .A1(n7105), .B0(n4404), .B1(n4170), .Y(n4574) );
  OAI22XL U3283 ( .A0(n4169), .A1(n7106), .B0(n4405), .B1(n4170), .Y(n4575) );
  OAI22XL U3284 ( .A0(n4169), .A1(n7107), .B0(n4406), .B1(n4170), .Y(n4576) );
  OAI22XL U3285 ( .A0(n4169), .A1(n7108), .B0(n4407), .B1(n4170), .Y(n4577) );
  OAI22XL U3286 ( .A0(n4169), .A1(n7109), .B0(n4408), .B1(n4171), .Y(n4578) );
  OAI22XL U3287 ( .A0(n1296), .A1(n7110), .B0(n4409), .B1(n6857), .Y(n4579) );
  OAI22XL U3288 ( .A0(n1296), .A1(n7111), .B0(n4410), .B1(n4170), .Y(n4580) );
  OAI22XL U3289 ( .A0(n4169), .A1(n7112), .B0(n4411), .B1(n4171), .Y(n4581) );
  OAI22XL U3290 ( .A0(n4169), .A1(n7113), .B0(n4412), .B1(n4171), .Y(n4582) );
  OAI22XL U3291 ( .A0(n4169), .A1(n7114), .B0(n4413), .B1(n4171), .Y(n4583) );
  OAI22XL U3292 ( .A0(n1296), .A1(n7115), .B0(n4414), .B1(n4170), .Y(n4584) );
  OAI22XL U3293 ( .A0(n4169), .A1(n7116), .B0(n4415), .B1(n4171), .Y(n4585) );
  OAI22XL U3294 ( .A0(n4169), .A1(n7117), .B0(n4416), .B1(n4171), .Y(n4586) );
  OAI22XL U3295 ( .A0(n4169), .A1(n7118), .B0(n4417), .B1(n4171), .Y(n4587) );
  OAI22XL U3296 ( .A0(n4169), .A1(n7119), .B0(n4418), .B1(n4171), .Y(n4588) );
  OAI22XL U3297 ( .A0(n4169), .A1(n7120), .B0(n4419), .B1(n4171), .Y(n4589) );
  OAI2BB2XL U3298 ( .B0(n4420), .B1(n4171), .A0N(n4170), .A1N(n1301), .Y(n4590) );
  OAI22XL U3299 ( .A0(n4172), .A1(n7072), .B0(n4396), .B1(n4173), .Y(n4591) );
  OAI22XL U3300 ( .A0(n4172), .A1(n7073), .B0(n4397), .B1(n4173), .Y(n4592) );
  OAI22XL U3301 ( .A0(n4172), .A1(n7074), .B0(n4398), .B1(n4173), .Y(n4593) );
  OAI22XL U3302 ( .A0(n4172), .A1(n7075), .B0(n4399), .B1(n4174), .Y(n4594) );
  OAI22XL U3303 ( .A0(n4172), .A1(n7076), .B0(n4400), .B1(n4174), .Y(n4595) );
  OAI22XL U3304 ( .A0(n4172), .A1(n7077), .B0(n4401), .B1(n4174), .Y(n4596) );
  OAI22XL U3305 ( .A0(n4172), .A1(n7078), .B0(n4402), .B1(n4173), .Y(n4597) );
  OAI22XL U3306 ( .A0(n4172), .A1(n7079), .B0(n4403), .B1(n6860), .Y(n4598) );
  OAI22XL U3307 ( .A0(n4172), .A1(n7080), .B0(n4404), .B1(n6860), .Y(n4599) );
  OAI22XL U3308 ( .A0(n4172), .A1(n7081), .B0(n4405), .B1(n4174), .Y(n4600) );
  OAI22XL U3309 ( .A0(n4172), .A1(n7082), .B0(n4406), .B1(n4173), .Y(n4601) );
  OAI22XL U3310 ( .A0(n4172), .A1(n7083), .B0(n4407), .B1(n4174), .Y(n4602) );
  OAI22XL U3311 ( .A0(n4172), .A1(n7084), .B0(n4408), .B1(n4174), .Y(n4603) );
  OAI22XL U3312 ( .A0(n4172), .A1(n7085), .B0(n4409), .B1(n4174), .Y(n4604) );
  OAI22XL U3313 ( .A0(n4172), .A1(n7086), .B0(n4410), .B1(n4174), .Y(n4605) );
  OAI22XL U3314 ( .A0(n4172), .A1(n7087), .B0(n4411), .B1(n4174), .Y(n4606) );
  OAI22XL U3315 ( .A0(n4172), .A1(n7088), .B0(n4412), .B1(n4174), .Y(n4607) );
  OAI22XL U3316 ( .A0(n4172), .A1(n7089), .B0(n4413), .B1(n4173), .Y(n4608) );
  OAI22XL U3317 ( .A0(n4172), .A1(n7090), .B0(n4414), .B1(n4173), .Y(n4609) );
  OAI22XL U3318 ( .A0(n4172), .A1(n7091), .B0(n4415), .B1(n4174), .Y(n4610) );
  OAI22XL U3319 ( .A0(n4172), .A1(n7092), .B0(n4416), .B1(n4173), .Y(n4611) );
  OAI22XL U3320 ( .A0(n1294), .A1(n7093), .B0(n4417), .B1(n4173), .Y(n4612) );
  OAI22XL U3321 ( .A0(n1294), .A1(n7094), .B0(n4418), .B1(n4173), .Y(n4613) );
  OAI22XL U3322 ( .A0(n1294), .A1(n7095), .B0(n4419), .B1(n4173), .Y(n4614) );
  OAI2BB2XL U3323 ( .B0(n4420), .B1(n4174), .A0N(n4173), .A1N(n1302), .Y(n4615) );
  OAI22XL U3324 ( .A0(n1295), .A1(n7047), .B0(n4396), .B1(n4176), .Y(n4422) );
  NAND2X1 U3325 ( .A(n8271), .B(n6831), .Y(n6843) );
  OAI21XL U3326 ( .A0(n4145), .A1(n6844), .B0(n8288), .Y(n4425) );
  OAI21XL U3327 ( .A0(n4135), .A1(n6844), .B0(n8287), .Y(n4426) );
  OAI21XL U3328 ( .A0(n4125), .A1(n6844), .B0(n8286), .Y(n4427) );
  OAI21XL U3329 ( .A0(n4115), .A1(n6844), .B0(n8285), .Y(n4428) );
  OAI21XL U3330 ( .A0(n1356), .A1(n6844), .B0(n8284), .Y(n4429) );
  OAI21XL U3331 ( .A0(n1697), .A1(n6844), .B0(n8283), .Y(n4430) );
  OAI21XL U3332 ( .A0(n1349), .A1(n6844), .B0(n8282), .Y(n4431) );
  OAI21XL U3333 ( .A0(n3998), .A1(n6844), .B0(n8281), .Y(n4432) );
  OAI21XL U3334 ( .A0(n3998), .A1(n1336), .B0(n8273), .Y(n4433) );
  OAI21XL U3335 ( .A0(n1697), .A1(n1336), .B0(n8275), .Y(n4435) );
  OAI21XL U3336 ( .A0(n1349), .A1(n1336), .B0(n8274), .Y(n4434) );
  OAI21XL U3337 ( .A0(n1355), .A1(n1336), .B0(n8276), .Y(n4436) );
  OAI21XL U3338 ( .A0(n4115), .A1(n1336), .B0(n8277), .Y(n4437) );
  OAI21XL U3339 ( .A0(n4135), .A1(n1336), .B0(n8279), .Y(n4439) );
  OAI21XL U3340 ( .A0(n4125), .A1(n1336), .B0(n8278), .Y(n4438) );
  OAI21XL U3341 ( .A0(n4145), .A1(n1336), .B0(n8280), .Y(n4440) );
  CLKINVX1 U3342 ( .A(mem_ready), .Y(n4421) );
  CLKBUFX3 U3343 ( .A(n6848), .Y(n1336) );
  NAND3X1 U3344 ( .A(n7045), .B(n8272), .C(n6839), .Y(n6848) );
  OAI2BB2XL U3345 ( .B0(n4420), .B1(n4162), .A0N(n4161), .A1N(n1303), .Y(n4515) );
  OAI2BB2XL U3346 ( .B0(n4420), .B1(n4165), .A0N(n4164), .A1N(n1304), .Y(n4540) );
  CLKINVX1 U3347 ( .A(proc_read), .Y(n4355) );
  NAND2X1 U3348 ( .A(proc_write), .B(n4355), .Y(n6831) );
  BUFX12 U3349 ( .A(proc_addr[3]), .Y(mem_addr[1]) );
  BUFX12 U3350 ( .A(proc_addr[2]), .Y(mem_addr[0]) );
endmodule


module CHIP ( clk, rst_n, mem_read_D, mem_write_D, mem_addr_D, mem_wdata_D, 
        mem_rdata_D, mem_ready_D, mem_read_I, mem_write_I, mem_addr_I, 
        mem_wdata_I, mem_rdata_I, mem_ready_I, DCACHE_addr, DCACHE_wdata, 
        DCACHE_wen );
  output [31:4] mem_addr_D;
  output [127:0] mem_wdata_D;
  input [127:0] mem_rdata_D;
  output [31:4] mem_addr_I;
  output [127:0] mem_wdata_I;
  input [127:0] mem_rdata_I;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input clk, rst_n, mem_ready_D, mem_ready_I;
  output mem_read_D, mem_write_D, mem_read_I, mem_write_I, DCACHE_wen;
  wire   ICACHE_stall, DCACHE_ren, DCACHE_stall, n2, n3;
  wire   [29:0] ICACHE_addr;
  wire   [31:0] ICACHE_wdata;
  wire   [31:0] ICACHE_rdata;
  wire   [31:0] DCACHE_rdata;

  MIPS_Pipeline i_MIPS ( .i_clk(clk), .rst_n(n2), .ICACHE_addr(ICACHE_addr), 
        .ICACHE_stall(ICACHE_stall), .ICACHE_rdata(ICACHE_rdata), .DCACHE_ren(
        DCACHE_ren), .DCACHE_wen(DCACHE_wen), .DCACHE_addr(DCACHE_addr), 
        .DCACHE_wdata(DCACHE_wdata), .DCACHE_stall(DCACHE_stall), 
        .DCACHE_rdata(DCACHE_rdata) );
  cache_0 D_cache ( .clk(clk), .proc_reset(n3), .proc_read(DCACHE_ren), 
        .proc_write(DCACHE_wen), .proc_addr(DCACHE_addr), .proc_wdata(
        DCACHE_wdata), .proc_stall(DCACHE_stall), .proc_rdata(DCACHE_rdata), 
        .mem_read(mem_read_D), .mem_write(mem_write_D), .mem_addr(mem_addr_D), 
        .mem_rdata(mem_rdata_D), .mem_wdata(mem_wdata_D), .mem_ready(
        mem_ready_D) );
  cache_1 I_cache ( .clk(clk), .proc_reset(n3), .proc_read(1'b1), .proc_write(
        1'b0), .proc_addr(ICACHE_addr), .proc_wdata({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .proc_stall(ICACHE_stall), .proc_rdata(
        ICACHE_rdata), .mem_read(mem_read_I), .mem_write(mem_write_I), 
        .mem_addr(mem_addr_I), .mem_rdata(mem_rdata_I), .mem_wdata(mem_wdata_I), .mem_ready(mem_ready_I) );
  CLKINVX1 U2 ( .A(n2), .Y(n3) );
  CLKBUFX3 U3 ( .A(rst_n), .Y(n2) );
endmodule

